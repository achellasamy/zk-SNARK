
module omega(wout);

    output [7:0] wout [0:63][0:63];

    assign wout[0][0] = 8'h00;
    assign wout[0][1] = 8'h00;
    assign wout[0][2] = 8'h00;
    assign wout[0][3] = 8'h00;
    assign wout[0][4] = 8'h00;
    assign wout[0][5] = 8'h00;
    assign wout[0][6] = 8'h00;
    assign wout[0][7] = 8'h00;
    assign wout[0][8] = 8'h00;
    assign wout[0][9] = 8'h00;
    assign wout[0][10] = 8'h00;
    assign wout[0][11] = 8'h00;
    assign wout[0][12] = 8'h00;
    assign wout[0][13] = 8'h00;
    assign wout[0][14] = 8'h00;
    assign wout[0][15] = 8'h00;
    assign wout[0][16] = 8'h00;
    assign wout[0][17] = 8'h00;
    assign wout[0][18] = 8'h00;
    assign wout[0][19] = 8'h00;
    assign wout[0][20] = 8'h00;
    assign wout[0][21] = 8'h00;
    assign wout[0][22] = 8'h00;
    assign wout[0][23] = 8'h00;
    assign wout[0][24] = 8'h00;
    assign wout[0][25] = 8'h00;
    assign wout[0][26] = 8'h00;
    assign wout[0][27] = 8'h00;
    assign wout[0][28] = 8'h00;
    assign wout[0][29] = 8'h00;
    assign wout[0][30] = 8'h00;
    assign wout[0][31] = 8'h00;
    assign wout[0][32] = 8'h00;
    assign wout[0][33] = 8'h00;
    assign wout[0][34] = 8'h00;
    assign wout[0][35] = 8'h00;
    assign wout[0][36] = 8'h00;
    assign wout[0][37] = 8'h00;
    assign wout[0][38] = 8'h00;
    assign wout[0][39] = 8'h00;
    assign wout[0][40] = 8'h00;
    assign wout[0][41] = 8'h00;
    assign wout[0][42] = 8'h00;
    assign wout[0][43] = 8'h00;
    assign wout[0][44] = 8'h00;
    assign wout[0][45] = 8'h00;
    assign wout[0][46] = 8'h00;
    assign wout[0][47] = 8'h00;
    assign wout[0][48] = 8'h00;
    assign wout[0][49] = 8'h00;
    assign wout[0][50] = 8'h00;
    assign wout[0][51] = 8'h00;
    assign wout[0][52] = 8'h00;
    assign wout[0][53] = 8'h00;
    assign wout[0][54] = 8'h00;
    assign wout[0][55] = 8'h00;
    assign wout[0][56] = 8'h00;
    assign wout[0][57] = 8'h00;
    assign wout[0][58] = 8'h00;
    assign wout[0][59] = 8'h00;
    assign wout[0][60] = 8'h00;
    assign wout[0][61] = 8'h00;
    assign wout[0][62] = 8'h00;
    assign wout[0][63] = 8'h00;
    assign wout[1][0] = 8'h00;
    assign wout[1][1] = 8'h01;
    assign wout[1][2] = 8'h02;
    assign wout[1][3] = 8'h03;
    assign wout[1][4] = 8'h04;
    assign wout[1][5] = 8'h05;
    assign wout[1][6] = 8'h06;
    assign wout[1][7] = 8'h07;
    assign wout[1][8] = 8'h08;
    assign wout[1][9] = 8'h09;
    assign wout[1][10] = 8'h0A;
    assign wout[1][11] = 8'h0B;
    assign wout[1][12] = 8'h0C;
    assign wout[1][13] = 8'h0D;
    assign wout[1][14] = 8'h0E;
    assign wout[1][15] = 8'h0F;
    assign wout[1][16] = 8'h10;
    assign wout[1][17] = 8'h11;
    assign wout[1][18] = 8'h12;
    assign wout[1][19] = 8'h13;
    assign wout[1][20] = 8'h14;
    assign wout[1][21] = 8'h15;
    assign wout[1][22] = 8'h16;
    assign wout[1][23] = 8'h17;
    assign wout[1][24] = 8'h18;
    assign wout[1][25] = 8'h19;
    assign wout[1][26] = 8'h1A;
    assign wout[1][27] = 8'h1B;
    assign wout[1][28] = 8'h1C;
    assign wout[1][29] = 8'h1D;
    assign wout[1][30] = 8'h1E;
    assign wout[1][31] = 8'h1F;
    assign wout[1][32] = 8'h20;
    assign wout[1][33] = 8'h21;
    assign wout[1][34] = 8'h22;
    assign wout[1][35] = 8'h23;
    assign wout[1][36] = 8'h24;
    assign wout[1][37] = 8'h25;
    assign wout[1][38] = 8'h26;
    assign wout[1][39] = 8'h27;
    assign wout[1][40] = 8'h28;
    assign wout[1][41] = 8'h29;
    assign wout[1][42] = 8'h2A;
    assign wout[1][43] = 8'h2B;
    assign wout[1][44] = 8'h2C;
    assign wout[1][45] = 8'h2D;
    assign wout[1][46] = 8'h2E;
    assign wout[1][47] = 8'h2F;
    assign wout[1][48] = 8'h30;
    assign wout[1][49] = 8'h31;
    assign wout[1][50] = 8'h32;
    assign wout[1][51] = 8'h33;
    assign wout[1][52] = 8'h34;
    assign wout[1][53] = 8'h35;
    assign wout[1][54] = 8'h36;
    assign wout[1][55] = 8'h37;
    assign wout[1][56] = 8'h38;
    assign wout[1][57] = 8'h39;
    assign wout[1][58] = 8'h3A;
    assign wout[1][59] = 8'h3B;
    assign wout[1][60] = 8'h3C;
    assign wout[1][61] = 8'h3D;
    assign wout[1][62] = 8'h3E;
    assign wout[1][63] = 8'h3F;
    assign wout[2][0] = 8'h00;
    assign wout[2][1] = 8'h02;
    assign wout[2][2] = 8'h04;
    assign wout[2][3] = 8'h06;
    assign wout[2][4] = 8'h08;
    assign wout[2][5] = 8'h0A;
    assign wout[2][6] = 8'h0C;
    assign wout[2][7] = 8'h0E;
    assign wout[2][8] = 8'h10;
    assign wout[2][9] = 8'h12;
    assign wout[2][10] = 8'h14;
    assign wout[2][11] = 8'h16;
    assign wout[2][12] = 8'h18;
    assign wout[2][13] = 8'h1A;
    assign wout[2][14] = 8'h1C;
    assign wout[2][15] = 8'h1E;
    assign wout[2][16] = 8'h20;
    assign wout[2][17] = 8'h22;
    assign wout[2][18] = 8'h24;
    assign wout[2][19] = 8'h26;
    assign wout[2][20] = 8'h28;
    assign wout[2][21] = 8'h2A;
    assign wout[2][22] = 8'h2C;
    assign wout[2][23] = 8'h2E;
    assign wout[2][24] = 8'h30;
    assign wout[2][25] = 8'h32;
    assign wout[2][26] = 8'h34;
    assign wout[2][27] = 8'h36;
    assign wout[2][28] = 8'h38;
    assign wout[2][29] = 8'h3A;
    assign wout[2][30] = 8'h3C;
    assign wout[2][31] = 8'h3E;
    assign wout[2][32] = 8'h40;
    assign wout[2][33] = 8'h42;
    assign wout[2][34] = 8'h44;
    assign wout[2][35] = 8'h46;
    assign wout[2][36] = 8'h48;
    assign wout[2][37] = 8'h4A;
    assign wout[2][38] = 8'h4C;
    assign wout[2][39] = 8'h4E;
    assign wout[2][40] = 8'h50;
    assign wout[2][41] = 8'h52;
    assign wout[2][42] = 8'h54;
    assign wout[2][43] = 8'h56;
    assign wout[2][44] = 8'h58;
    assign wout[2][45] = 8'h5A;
    assign wout[2][46] = 8'h5C;
    assign wout[2][47] = 8'h5E;
    assign wout[2][48] = 8'h60;
    assign wout[2][49] = 8'h62;
    assign wout[2][50] = 8'h64;
    assign wout[2][51] = 8'h66;
    assign wout[2][52] = 8'h68;
    assign wout[2][53] = 8'h6A;
    assign wout[2][54] = 8'h6C;
    assign wout[2][55] = 8'h6E;
    assign wout[2][56] = 8'h70;
    assign wout[2][57] = 8'h72;
    assign wout[2][58] = 8'h74;
    assign wout[2][59] = 8'h76;
    assign wout[2][60] = 8'h78;
    assign wout[2][61] = 8'h7A;
    assign wout[2][62] = 8'h7C;
    assign wout[2][63] = 8'h7E;
    assign wout[3][0] = 8'h00;
    assign wout[3][1] = 8'h03;
    assign wout[3][2] = 8'h06;
    assign wout[3][3] = 8'h09;
    assign wout[3][4] = 8'h0C;
    assign wout[3][5] = 8'h0F;
    assign wout[3][6] = 8'h12;
    assign wout[3][7] = 8'h15;
    assign wout[3][8] = 8'h18;
    assign wout[3][9] = 8'h1B;
    assign wout[3][10] = 8'h1E;
    assign wout[3][11] = 8'h21;
    assign wout[3][12] = 8'h24;
    assign wout[3][13] = 8'h27;
    assign wout[3][14] = 8'h2A;
    assign wout[3][15] = 8'h2D;
    assign wout[3][16] = 8'h30;
    assign wout[3][17] = 8'h33;
    assign wout[3][18] = 8'h36;
    assign wout[3][19] = 8'h39;
    assign wout[3][20] = 8'h3C;
    assign wout[3][21] = 8'h3F;
    assign wout[3][22] = 8'h42;
    assign wout[3][23] = 8'h45;
    assign wout[3][24] = 8'h48;
    assign wout[3][25] = 8'h4B;
    assign wout[3][26] = 8'h4E;
    assign wout[3][27] = 8'h51;
    assign wout[3][28] = 8'h54;
    assign wout[3][29] = 8'h57;
    assign wout[3][30] = 8'h5A;
    assign wout[3][31] = 8'h5D;
    assign wout[3][32] = 8'h60;
    assign wout[3][33] = 8'h63;
    assign wout[3][34] = 8'h66;
    assign wout[3][35] = 8'h69;
    assign wout[3][36] = 8'h6C;
    assign wout[3][37] = 8'h6F;
    assign wout[3][38] = 8'h72;
    assign wout[3][39] = 8'h75;
    assign wout[3][40] = 8'h78;
    assign wout[3][41] = 8'h7B;
    assign wout[3][42] = 8'h7E;
    assign wout[3][43] = 8'h81;
    assign wout[3][44] = 8'h84;
    assign wout[3][45] = 8'h87;
    assign wout[3][46] = 8'h8A;
    assign wout[3][47] = 8'h8D;
    assign wout[3][48] = 8'h90;
    assign wout[3][49] = 8'h93;
    assign wout[3][50] = 8'h96;
    assign wout[3][51] = 8'h99;
    assign wout[3][52] = 8'h9C;
    assign wout[3][53] = 8'h9F;
    assign wout[3][54] = 8'hA2;
    assign wout[3][55] = 8'hA5;
    assign wout[3][56] = 8'hA8;
    assign wout[3][57] = 8'hAB;
    assign wout[3][58] = 8'hAE;
    assign wout[3][59] = 8'hB1;
    assign wout[3][60] = 8'hB4;
    assign wout[3][61] = 8'hB7;
    assign wout[3][62] = 8'hBA;
    assign wout[3][63] = 8'hBD;
    assign wout[4][0] = 8'h00;
    assign wout[4][1] = 8'h04;
    assign wout[4][2] = 8'h08;
    assign wout[4][3] = 8'h0C;
    assign wout[4][4] = 8'h10;
    assign wout[4][5] = 8'h14;
    assign wout[4][6] = 8'h18;
    assign wout[4][7] = 8'h1C;
    assign wout[4][8] = 8'h20;
    assign wout[4][9] = 8'h24;
    assign wout[4][10] = 8'h28;
    assign wout[4][11] = 8'h2C;
    assign wout[4][12] = 8'h30;
    assign wout[4][13] = 8'h34;
    assign wout[4][14] = 8'h38;
    assign wout[4][15] = 8'h3C;
    assign wout[4][16] = 8'h40;
    assign wout[4][17] = 8'h44;
    assign wout[4][18] = 8'h48;
    assign wout[4][19] = 8'h4C;
    assign wout[4][20] = 8'h50;
    assign wout[4][21] = 8'h54;
    assign wout[4][22] = 8'h58;
    assign wout[4][23] = 8'h5C;
    assign wout[4][24] = 8'h60;
    assign wout[4][25] = 8'h64;
    assign wout[4][26] = 8'h68;
    assign wout[4][27] = 8'h6C;
    assign wout[4][28] = 8'h70;
    assign wout[4][29] = 8'h74;
    assign wout[4][30] = 8'h78;
    assign wout[4][31] = 8'h7C;
    assign wout[4][32] = 8'h80;
    assign wout[4][33] = 8'h84;
    assign wout[4][34] = 8'h88;
    assign wout[4][35] = 8'h8C;
    assign wout[4][36] = 8'h90;
    assign wout[4][37] = 8'h94;
    assign wout[4][38] = 8'h98;
    assign wout[4][39] = 8'h9C;
    assign wout[4][40] = 8'hA0;
    assign wout[4][41] = 8'hA4;
    assign wout[4][42] = 8'hA8;
    assign wout[4][43] = 8'hAC;
    assign wout[4][44] = 8'hB0;
    assign wout[4][45] = 8'hB4;
    assign wout[4][46] = 8'hB8;
    assign wout[4][47] = 8'hBC;
    assign wout[4][48] = 8'hC0;
    assign wout[4][49] = 8'hC4;
    assign wout[4][50] = 8'hC8;
    assign wout[4][51] = 8'hCC;
    assign wout[4][52] = 8'hD0;
    assign wout[4][53] = 8'hD4;
    assign wout[4][54] = 8'hD8;
    assign wout[4][55] = 8'hDC;
    assign wout[4][56] = 8'hE0;
    assign wout[4][57] = 8'hE4;
    assign wout[4][58] = 8'hE8;
    assign wout[4][59] = 8'hEC;
    assign wout[4][60] = 8'hF0;
    assign wout[4][61] = 8'hF4;
    assign wout[4][62] = 8'hF8;
    assign wout[4][63] = 8'hFC;
    assign wout[5][0] = 8'h00;
    assign wout[5][1] = 8'h05;
    assign wout[5][2] = 8'h0A;
    assign wout[5][3] = 8'h0F;
    assign wout[5][4] = 8'h14;
    assign wout[5][5] = 8'h19;
    assign wout[5][6] = 8'h1E;
    assign wout[5][7] = 8'h23;
    assign wout[5][8] = 8'h28;
    assign wout[5][9] = 8'h2D;
    assign wout[5][10] = 8'h32;
    assign wout[5][11] = 8'h37;
    assign wout[5][12] = 8'h3C;
    assign wout[5][13] = 8'h41;
    assign wout[5][14] = 8'h46;
    assign wout[5][15] = 8'h4B;
    assign wout[5][16] = 8'h50;
    assign wout[5][17] = 8'h55;
    assign wout[5][18] = 8'h5A;
    assign wout[5][19] = 8'h5F;
    assign wout[5][20] = 8'h64;
    assign wout[5][21] = 8'h69;
    assign wout[5][22] = 8'h6E;
    assign wout[5][23] = 8'h73;
    assign wout[5][24] = 8'h78;
    assign wout[5][25] = 8'h7D;
    assign wout[5][26] = 8'h82;
    assign wout[5][27] = 8'h87;
    assign wout[5][28] = 8'h8C;
    assign wout[5][29] = 8'h91;
    assign wout[5][30] = 8'h96;
    assign wout[5][31] = 8'h9B;
    assign wout[5][32] = 8'hA0;
    assign wout[5][33] = 8'hA5;
    assign wout[5][34] = 8'hAA;
    assign wout[5][35] = 8'hAF;
    assign wout[5][36] = 8'hB4;
    assign wout[5][37] = 8'hB9;
    assign wout[5][38] = 8'hBE;
    assign wout[5][39] = 8'hC3;
    assign wout[5][40] = 8'hC8;
    assign wout[5][41] = 8'hCD;
    assign wout[5][42] = 8'hD2;
    assign wout[5][43] = 8'hD7;
    assign wout[5][44] = 8'hDC;
    assign wout[5][45] = 8'hE1;
    assign wout[5][46] = 8'hE6;
    assign wout[5][47] = 8'hEB;
    assign wout[5][48] = 8'hF0;
    assign wout[5][49] = 8'hF5;
    assign wout[5][50] = 8'hFA;
    assign wout[5][51] = 8'hFF;
    assign wout[5][52] = 8'h04;
    assign wout[5][53] = 8'h09;
    assign wout[5][54] = 8'h0E;
    assign wout[5][55] = 8'h13;
    assign wout[5][56] = 8'h18;
    assign wout[5][57] = 8'h1D;
    assign wout[5][58] = 8'h22;
    assign wout[5][59] = 8'h27;
    assign wout[5][60] = 8'h2C;
    assign wout[5][61] = 8'h31;
    assign wout[5][62] = 8'h36;
    assign wout[5][63] = 8'h3B;
    assign wout[6][0] = 8'h00;
    assign wout[6][1] = 8'h06;
    assign wout[6][2] = 8'h0C;
    assign wout[6][3] = 8'h12;
    assign wout[6][4] = 8'h18;
    assign wout[6][5] = 8'h1E;
    assign wout[6][6] = 8'h24;
    assign wout[6][7] = 8'h2A;
    assign wout[6][8] = 8'h30;
    assign wout[6][9] = 8'h36;
    assign wout[6][10] = 8'h3C;
    assign wout[6][11] = 8'h42;
    assign wout[6][12] = 8'h48;
    assign wout[6][13] = 8'h4E;
    assign wout[6][14] = 8'h54;
    assign wout[6][15] = 8'h5A;
    assign wout[6][16] = 8'h60;
    assign wout[6][17] = 8'h66;
    assign wout[6][18] = 8'h6C;
    assign wout[6][19] = 8'h72;
    assign wout[6][20] = 8'h78;
    assign wout[6][21] = 8'h7E;
    assign wout[6][22] = 8'h84;
    assign wout[6][23] = 8'h8A;
    assign wout[6][24] = 8'h90;
    assign wout[6][25] = 8'h96;
    assign wout[6][26] = 8'h9C;
    assign wout[6][27] = 8'hA2;
    assign wout[6][28] = 8'hA8;
    assign wout[6][29] = 8'hAE;
    assign wout[6][30] = 8'hB4;
    assign wout[6][31] = 8'hBA;
    assign wout[6][32] = 8'hC0;
    assign wout[6][33] = 8'hC6;
    assign wout[6][34] = 8'hCC;
    assign wout[6][35] = 8'hD2;
    assign wout[6][36] = 8'hD8;
    assign wout[6][37] = 8'hDE;
    assign wout[6][38] = 8'hE4;
    assign wout[6][39] = 8'hEA;
    assign wout[6][40] = 8'hF0;
    assign wout[6][41] = 8'hF6;
    assign wout[6][42] = 8'hFC;
    assign wout[6][43] = 8'h02;
    assign wout[6][44] = 8'h08;
    assign wout[6][45] = 8'h0E;
    assign wout[6][46] = 8'h14;
    assign wout[6][47] = 8'h1A;
    assign wout[6][48] = 8'h20;
    assign wout[6][49] = 8'h26;
    assign wout[6][50] = 8'h2C;
    assign wout[6][51] = 8'h32;
    assign wout[6][52] = 8'h38;
    assign wout[6][53] = 8'h3E;
    assign wout[6][54] = 8'h44;
    assign wout[6][55] = 8'h4A;
    assign wout[6][56] = 8'h50;
    assign wout[6][57] = 8'h56;
    assign wout[6][58] = 8'h5C;
    assign wout[6][59] = 8'h62;
    assign wout[6][60] = 8'h68;
    assign wout[6][61] = 8'h6E;
    assign wout[6][62] = 8'h74;
    assign wout[6][63] = 8'h7A;
    assign wout[7][0] = 8'h00;
    assign wout[7][1] = 8'h07;
    assign wout[7][2] = 8'h0E;
    assign wout[7][3] = 8'h15;
    assign wout[7][4] = 8'h1C;
    assign wout[7][5] = 8'h23;
    assign wout[7][6] = 8'h2A;
    assign wout[7][7] = 8'h31;
    assign wout[7][8] = 8'h38;
    assign wout[7][9] = 8'h3F;
    assign wout[7][10] = 8'h46;
    assign wout[7][11] = 8'h4D;
    assign wout[7][12] = 8'h54;
    assign wout[7][13] = 8'h5B;
    assign wout[7][14] = 8'h62;
    assign wout[7][15] = 8'h69;
    assign wout[7][16] = 8'h70;
    assign wout[7][17] = 8'h77;
    assign wout[7][18] = 8'h7E;
    assign wout[7][19] = 8'h85;
    assign wout[7][20] = 8'h8C;
    assign wout[7][21] = 8'h93;
    assign wout[7][22] = 8'h9A;
    assign wout[7][23] = 8'hA1;
    assign wout[7][24] = 8'hA8;
    assign wout[7][25] = 8'hAF;
    assign wout[7][26] = 8'hB6;
    assign wout[7][27] = 8'hBD;
    assign wout[7][28] = 8'hC4;
    assign wout[7][29] = 8'hCB;
    assign wout[7][30] = 8'hD2;
    assign wout[7][31] = 8'hD9;
    assign wout[7][32] = 8'hE0;
    assign wout[7][33] = 8'hE7;
    assign wout[7][34] = 8'hEE;
    assign wout[7][35] = 8'hF5;
    assign wout[7][36] = 8'hFC;
    assign wout[7][37] = 8'h03;
    assign wout[7][38] = 8'h0A;
    assign wout[7][39] = 8'h11;
    assign wout[7][40] = 8'h18;
    assign wout[7][41] = 8'h1F;
    assign wout[7][42] = 8'h26;
    assign wout[7][43] = 8'h2D;
    assign wout[7][44] = 8'h34;
    assign wout[7][45] = 8'h3B;
    assign wout[7][46] = 8'h42;
    assign wout[7][47] = 8'h49;
    assign wout[7][48] = 8'h50;
    assign wout[7][49] = 8'h57;
    assign wout[7][50] = 8'h5E;
    assign wout[7][51] = 8'h65;
    assign wout[7][52] = 8'h6C;
    assign wout[7][53] = 8'h73;
    assign wout[7][54] = 8'h7A;
    assign wout[7][55] = 8'h81;
    assign wout[7][56] = 8'h88;
    assign wout[7][57] = 8'h8F;
    assign wout[7][58] = 8'h96;
    assign wout[7][59] = 8'h9D;
    assign wout[7][60] = 8'hA4;
    assign wout[7][61] = 8'hAB;
    assign wout[7][62] = 8'hB2;
    assign wout[7][63] = 8'hB9;
    assign wout[8][0] = 8'h00;
    assign wout[8][1] = 8'h08;
    assign wout[8][2] = 8'h10;
    assign wout[8][3] = 8'h18;
    assign wout[8][4] = 8'h20;
    assign wout[8][5] = 8'h28;
    assign wout[8][6] = 8'h30;
    assign wout[8][7] = 8'h38;
    assign wout[8][8] = 8'h40;
    assign wout[8][9] = 8'h48;
    assign wout[8][10] = 8'h50;
    assign wout[8][11] = 8'h58;
    assign wout[8][12] = 8'h60;
    assign wout[8][13] = 8'h68;
    assign wout[8][14] = 8'h70;
    assign wout[8][15] = 8'h78;
    assign wout[8][16] = 8'h80;
    assign wout[8][17] = 8'h88;
    assign wout[8][18] = 8'h90;
    assign wout[8][19] = 8'h98;
    assign wout[8][20] = 8'hA0;
    assign wout[8][21] = 8'hA8;
    assign wout[8][22] = 8'hB0;
    assign wout[8][23] = 8'hB8;
    assign wout[8][24] = 8'hC0;
    assign wout[8][25] = 8'hC8;
    assign wout[8][26] = 8'hD0;
    assign wout[8][27] = 8'hD8;
    assign wout[8][28] = 8'hE0;
    assign wout[8][29] = 8'hE8;
    assign wout[8][30] = 8'hF0;
    assign wout[8][31] = 8'hF8;
    assign wout[8][32] = 8'h00;
    assign wout[8][33] = 8'h08;
    assign wout[8][34] = 8'h10;
    assign wout[8][35] = 8'h18;
    assign wout[8][36] = 8'h20;
    assign wout[8][37] = 8'h28;
    assign wout[8][38] = 8'h30;
    assign wout[8][39] = 8'h38;
    assign wout[8][40] = 8'h40;
    assign wout[8][41] = 8'h48;
    assign wout[8][42] = 8'h50;
    assign wout[8][43] = 8'h58;
    assign wout[8][44] = 8'h60;
    assign wout[8][45] = 8'h68;
    assign wout[8][46] = 8'h70;
    assign wout[8][47] = 8'h78;
    assign wout[8][48] = 8'h80;
    assign wout[8][49] = 8'h88;
    assign wout[8][50] = 8'h90;
    assign wout[8][51] = 8'h98;
    assign wout[8][52] = 8'hA0;
    assign wout[8][53] = 8'hA8;
    assign wout[8][54] = 8'hB0;
    assign wout[8][55] = 8'hB8;
    assign wout[8][56] = 8'hC0;
    assign wout[8][57] = 8'hC8;
    assign wout[8][58] = 8'hD0;
    assign wout[8][59] = 8'hD8;
    assign wout[8][60] = 8'hE0;
    assign wout[8][61] = 8'hE8;
    assign wout[8][62] = 8'hF0;
    assign wout[8][63] = 8'hF8;
    assign wout[9][0] = 8'h00;
    assign wout[9][1] = 8'h09;
    assign wout[9][2] = 8'h12;
    assign wout[9][3] = 8'h1B;
    assign wout[9][4] = 8'h24;
    assign wout[9][5] = 8'h2D;
    assign wout[9][6] = 8'h36;
    assign wout[9][7] = 8'h3F;
    assign wout[9][8] = 8'h48;
    assign wout[9][9] = 8'h51;
    assign wout[9][10] = 8'h5A;
    assign wout[9][11] = 8'h63;
    assign wout[9][12] = 8'h6C;
    assign wout[9][13] = 8'h75;
    assign wout[9][14] = 8'h7E;
    assign wout[9][15] = 8'h87;
    assign wout[9][16] = 8'h90;
    assign wout[9][17] = 8'h99;
    assign wout[9][18] = 8'hA2;
    assign wout[9][19] = 8'hAB;
    assign wout[9][20] = 8'hB4;
    assign wout[9][21] = 8'hBD;
    assign wout[9][22] = 8'hC6;
    assign wout[9][23] = 8'hCF;
    assign wout[9][24] = 8'hD8;
    assign wout[9][25] = 8'hE1;
    assign wout[9][26] = 8'hEA;
    assign wout[9][27] = 8'hF3;
    assign wout[9][28] = 8'hFC;
    assign wout[9][29] = 8'h05;
    assign wout[9][30] = 8'h0E;
    assign wout[9][31] = 8'h17;
    assign wout[9][32] = 8'h20;
    assign wout[9][33] = 8'h29;
    assign wout[9][34] = 8'h32;
    assign wout[9][35] = 8'h3B;
    assign wout[9][36] = 8'h44;
    assign wout[9][37] = 8'h4D;
    assign wout[9][38] = 8'h56;
    assign wout[9][39] = 8'h5F;
    assign wout[9][40] = 8'h68;
    assign wout[9][41] = 8'h71;
    assign wout[9][42] = 8'h7A;
    assign wout[9][43] = 8'h83;
    assign wout[9][44] = 8'h8C;
    assign wout[9][45] = 8'h95;
    assign wout[9][46] = 8'h9E;
    assign wout[9][47] = 8'hA7;
    assign wout[9][48] = 8'hB0;
    assign wout[9][49] = 8'hB9;
    assign wout[9][50] = 8'hC2;
    assign wout[9][51] = 8'hCB;
    assign wout[9][52] = 8'hD4;
    assign wout[9][53] = 8'hDD;
    assign wout[9][54] = 8'hE6;
    assign wout[9][55] = 8'hEF;
    assign wout[9][56] = 8'hF8;
    assign wout[9][57] = 8'h01;
    assign wout[9][58] = 8'h0A;
    assign wout[9][59] = 8'h13;
    assign wout[9][60] = 8'h1C;
    assign wout[9][61] = 8'h25;
    assign wout[9][62] = 8'h2E;
    assign wout[9][63] = 8'h37;
    assign wout[10][0] = 8'h00;
    assign wout[10][1] = 8'h0A;
    assign wout[10][2] = 8'h14;
    assign wout[10][3] = 8'h1E;
    assign wout[10][4] = 8'h28;
    assign wout[10][5] = 8'h32;
    assign wout[10][6] = 8'h3C;
    assign wout[10][7] = 8'h46;
    assign wout[10][8] = 8'h50;
    assign wout[10][9] = 8'h5A;
    assign wout[10][10] = 8'h64;
    assign wout[10][11] = 8'h6E;
    assign wout[10][12] = 8'h78;
    assign wout[10][13] = 8'h82;
    assign wout[10][14] = 8'h8C;
    assign wout[10][15] = 8'h96;
    assign wout[10][16] = 8'hA0;
    assign wout[10][17] = 8'hAA;
    assign wout[10][18] = 8'hB4;
    assign wout[10][19] = 8'hBE;
    assign wout[10][20] = 8'hC8;
    assign wout[10][21] = 8'hD2;
    assign wout[10][22] = 8'hDC;
    assign wout[10][23] = 8'hE6;
    assign wout[10][24] = 8'hF0;
    assign wout[10][25] = 8'hFA;
    assign wout[10][26] = 8'h04;
    assign wout[10][27] = 8'h0E;
    assign wout[10][28] = 8'h18;
    assign wout[10][29] = 8'h22;
    assign wout[10][30] = 8'h2C;
    assign wout[10][31] = 8'h36;
    assign wout[10][32] = 8'h40;
    assign wout[10][33] = 8'h4A;
    assign wout[10][34] = 8'h54;
    assign wout[10][35] = 8'h5E;
    assign wout[10][36] = 8'h68;
    assign wout[10][37] = 8'h72;
    assign wout[10][38] = 8'h7C;
    assign wout[10][39] = 8'h86;
    assign wout[10][40] = 8'h90;
    assign wout[10][41] = 8'h9A;
    assign wout[10][42] = 8'hA4;
    assign wout[10][43] = 8'hAE;
    assign wout[10][44] = 8'hB8;
    assign wout[10][45] = 8'hC2;
    assign wout[10][46] = 8'hCC;
    assign wout[10][47] = 8'hD6;
    assign wout[10][48] = 8'hE0;
    assign wout[10][49] = 8'hEA;
    assign wout[10][50] = 8'hF4;
    assign wout[10][51] = 8'hFE;
    assign wout[10][52] = 8'h08;
    assign wout[10][53] = 8'h12;
    assign wout[10][54] = 8'h1C;
    assign wout[10][55] = 8'h26;
    assign wout[10][56] = 8'h30;
    assign wout[10][57] = 8'h3A;
    assign wout[10][58] = 8'h44;
    assign wout[10][59] = 8'h4E;
    assign wout[10][60] = 8'h58;
    assign wout[10][61] = 8'h62;
    assign wout[10][62] = 8'h6C;
    assign wout[10][63] = 8'h76;
    assign wout[11][0] = 8'h00;
    assign wout[11][1] = 8'h0B;
    assign wout[11][2] = 8'h16;
    assign wout[11][3] = 8'h21;
    assign wout[11][4] = 8'h2C;
    assign wout[11][5] = 8'h37;
    assign wout[11][6] = 8'h42;
    assign wout[11][7] = 8'h4D;
    assign wout[11][8] = 8'h58;
    assign wout[11][9] = 8'h63;
    assign wout[11][10] = 8'h6E;
    assign wout[11][11] = 8'h79;
    assign wout[11][12] = 8'h84;
    assign wout[11][13] = 8'h8F;
    assign wout[11][14] = 8'h9A;
    assign wout[11][15] = 8'hA5;
    assign wout[11][16] = 8'hB0;
    assign wout[11][17] = 8'hBB;
    assign wout[11][18] = 8'hC6;
    assign wout[11][19] = 8'hD1;
    assign wout[11][20] = 8'hDC;
    assign wout[11][21] = 8'hE7;
    assign wout[11][22] = 8'hF2;
    assign wout[11][23] = 8'hFD;
    assign wout[11][24] = 8'h08;
    assign wout[11][25] = 8'h13;
    assign wout[11][26] = 8'h1E;
    assign wout[11][27] = 8'h29;
    assign wout[11][28] = 8'h34;
    assign wout[11][29] = 8'h3F;
    assign wout[11][30] = 8'h4A;
    assign wout[11][31] = 8'h55;
    assign wout[11][32] = 8'h60;
    assign wout[11][33] = 8'h6B;
    assign wout[11][34] = 8'h76;
    assign wout[11][35] = 8'h81;
    assign wout[11][36] = 8'h8C;
    assign wout[11][37] = 8'h97;
    assign wout[11][38] = 8'hA2;
    assign wout[11][39] = 8'hAD;
    assign wout[11][40] = 8'hB8;
    assign wout[11][41] = 8'hC3;
    assign wout[11][42] = 8'hCE;
    assign wout[11][43] = 8'hD9;
    assign wout[11][44] = 8'hE4;
    assign wout[11][45] = 8'hEF;
    assign wout[11][46] = 8'hFA;
    assign wout[11][47] = 8'h05;
    assign wout[11][48] = 8'h10;
    assign wout[11][49] = 8'h1B;
    assign wout[11][50] = 8'h26;
    assign wout[11][51] = 8'h31;
    assign wout[11][52] = 8'h3C;
    assign wout[11][53] = 8'h47;
    assign wout[11][54] = 8'h52;
    assign wout[11][55] = 8'h5D;
    assign wout[11][56] = 8'h68;
    assign wout[11][57] = 8'h73;
    assign wout[11][58] = 8'h7E;
    assign wout[11][59] = 8'h89;
    assign wout[11][60] = 8'h94;
    assign wout[11][61] = 8'h9F;
    assign wout[11][62] = 8'hAA;
    assign wout[11][63] = 8'hB5;
    assign wout[12][0] = 8'h00;
    assign wout[12][1] = 8'h0C;
    assign wout[12][2] = 8'h18;
    assign wout[12][3] = 8'h24;
    assign wout[12][4] = 8'h30;
    assign wout[12][5] = 8'h3C;
    assign wout[12][6] = 8'h48;
    assign wout[12][7] = 8'h54;
    assign wout[12][8] = 8'h60;
    assign wout[12][9] = 8'h6C;
    assign wout[12][10] = 8'h78;
    assign wout[12][11] = 8'h84;
    assign wout[12][12] = 8'h90;
    assign wout[12][13] = 8'h9C;
    assign wout[12][14] = 8'hA8;
    assign wout[12][15] = 8'hB4;
    assign wout[12][16] = 8'hC0;
    assign wout[12][17] = 8'hCC;
    assign wout[12][18] = 8'hD8;
    assign wout[12][19] = 8'hE4;
    assign wout[12][20] = 8'hF0;
    assign wout[12][21] = 8'hFC;
    assign wout[12][22] = 8'h08;
    assign wout[12][23] = 8'h14;
    assign wout[12][24] = 8'h20;
    assign wout[12][25] = 8'h2C;
    assign wout[12][26] = 8'h38;
    assign wout[12][27] = 8'h44;
    assign wout[12][28] = 8'h50;
    assign wout[12][29] = 8'h5C;
    assign wout[12][30] = 8'h68;
    assign wout[12][31] = 8'h74;
    assign wout[12][32] = 8'h80;
    assign wout[12][33] = 8'h8C;
    assign wout[12][34] = 8'h98;
    assign wout[12][35] = 8'hA4;
    assign wout[12][36] = 8'hB0;
    assign wout[12][37] = 8'hBC;
    assign wout[12][38] = 8'hC8;
    assign wout[12][39] = 8'hD4;
    assign wout[12][40] = 8'hE0;
    assign wout[12][41] = 8'hEC;
    assign wout[12][42] = 8'hF8;
    assign wout[12][43] = 8'h04;
    assign wout[12][44] = 8'h10;
    assign wout[12][45] = 8'h1C;
    assign wout[12][46] = 8'h28;
    assign wout[12][47] = 8'h34;
    assign wout[12][48] = 8'h40;
    assign wout[12][49] = 8'h4C;
    assign wout[12][50] = 8'h58;
    assign wout[12][51] = 8'h64;
    assign wout[12][52] = 8'h70;
    assign wout[12][53] = 8'h7C;
    assign wout[12][54] = 8'h88;
    assign wout[12][55] = 8'h94;
    assign wout[12][56] = 8'hA0;
    assign wout[12][57] = 8'hAC;
    assign wout[12][58] = 8'hB8;
    assign wout[12][59] = 8'hC4;
    assign wout[12][60] = 8'hD0;
    assign wout[12][61] = 8'hDC;
    assign wout[12][62] = 8'hE8;
    assign wout[12][63] = 8'hF4;
    assign wout[13][0] = 8'h00;
    assign wout[13][1] = 8'h0D;
    assign wout[13][2] = 8'h1A;
    assign wout[13][3] = 8'h27;
    assign wout[13][4] = 8'h34;
    assign wout[13][5] = 8'h41;
    assign wout[13][6] = 8'h4E;
    assign wout[13][7] = 8'h5B;
    assign wout[13][8] = 8'h68;
    assign wout[13][9] = 8'h75;
    assign wout[13][10] = 8'h82;
    assign wout[13][11] = 8'h8F;
    assign wout[13][12] = 8'h9C;
    assign wout[13][13] = 8'hA9;
    assign wout[13][14] = 8'hB6;
    assign wout[13][15] = 8'hC3;
    assign wout[13][16] = 8'hD0;
    assign wout[13][17] = 8'hDD;
    assign wout[13][18] = 8'hEA;
    assign wout[13][19] = 8'hF7;
    assign wout[13][20] = 8'h04;
    assign wout[13][21] = 8'h11;
    assign wout[13][22] = 8'h1E;
    assign wout[13][23] = 8'h2B;
    assign wout[13][24] = 8'h38;
    assign wout[13][25] = 8'h45;
    assign wout[13][26] = 8'h52;
    assign wout[13][27] = 8'h5F;
    assign wout[13][28] = 8'h6C;
    assign wout[13][29] = 8'h79;
    assign wout[13][30] = 8'h86;
    assign wout[13][31] = 8'h93;
    assign wout[13][32] = 8'hA0;
    assign wout[13][33] = 8'hAD;
    assign wout[13][34] = 8'hBA;
    assign wout[13][35] = 8'hC7;
    assign wout[13][36] = 8'hD4;
    assign wout[13][37] = 8'hE1;
    assign wout[13][38] = 8'hEE;
    assign wout[13][39] = 8'hFB;
    assign wout[13][40] = 8'h08;
    assign wout[13][41] = 8'h15;
    assign wout[13][42] = 8'h22;
    assign wout[13][43] = 8'h2F;
    assign wout[13][44] = 8'h3C;
    assign wout[13][45] = 8'h49;
    assign wout[13][46] = 8'h56;
    assign wout[13][47] = 8'h63;
    assign wout[13][48] = 8'h70;
    assign wout[13][49] = 8'h7D;
    assign wout[13][50] = 8'h8A;
    assign wout[13][51] = 8'h97;
    assign wout[13][52] = 8'hA4;
    assign wout[13][53] = 8'hB1;
    assign wout[13][54] = 8'hBE;
    assign wout[13][55] = 8'hCB;
    assign wout[13][56] = 8'hD8;
    assign wout[13][57] = 8'hE5;
    assign wout[13][58] = 8'hF2;
    assign wout[13][59] = 8'hFF;
    assign wout[13][60] = 8'h0C;
    assign wout[13][61] = 8'h19;
    assign wout[13][62] = 8'h26;
    assign wout[13][63] = 8'h33;
    assign wout[14][0] = 8'h00;
    assign wout[14][1] = 8'h0E;
    assign wout[14][2] = 8'h1C;
    assign wout[14][3] = 8'h2A;
    assign wout[14][4] = 8'h38;
    assign wout[14][5] = 8'h46;
    assign wout[14][6] = 8'h54;
    assign wout[14][7] = 8'h62;
    assign wout[14][8] = 8'h70;
    assign wout[14][9] = 8'h7E;
    assign wout[14][10] = 8'h8C;
    assign wout[14][11] = 8'h9A;
    assign wout[14][12] = 8'hA8;
    assign wout[14][13] = 8'hB6;
    assign wout[14][14] = 8'hC4;
    assign wout[14][15] = 8'hD2;
    assign wout[14][16] = 8'hE0;
    assign wout[14][17] = 8'hEE;
    assign wout[14][18] = 8'hFC;
    assign wout[14][19] = 8'h0A;
    assign wout[14][20] = 8'h18;
    assign wout[14][21] = 8'h26;
    assign wout[14][22] = 8'h34;
    assign wout[14][23] = 8'h42;
    assign wout[14][24] = 8'h50;
    assign wout[14][25] = 8'h5E;
    assign wout[14][26] = 8'h6C;
    assign wout[14][27] = 8'h7A;
    assign wout[14][28] = 8'h88;
    assign wout[14][29] = 8'h96;
    assign wout[14][30] = 8'hA4;
    assign wout[14][31] = 8'hB2;
    assign wout[14][32] = 8'hC0;
    assign wout[14][33] = 8'hCE;
    assign wout[14][34] = 8'hDC;
    assign wout[14][35] = 8'hEA;
    assign wout[14][36] = 8'hF8;
    assign wout[14][37] = 8'h06;
    assign wout[14][38] = 8'h14;
    assign wout[14][39] = 8'h22;
    assign wout[14][40] = 8'h30;
    assign wout[14][41] = 8'h3E;
    assign wout[14][42] = 8'h4C;
    assign wout[14][43] = 8'h5A;
    assign wout[14][44] = 8'h68;
    assign wout[14][45] = 8'h76;
    assign wout[14][46] = 8'h84;
    assign wout[14][47] = 8'h92;
    assign wout[14][48] = 8'hA0;
    assign wout[14][49] = 8'hAE;
    assign wout[14][50] = 8'hBC;
    assign wout[14][51] = 8'hCA;
    assign wout[14][52] = 8'hD8;
    assign wout[14][53] = 8'hE6;
    assign wout[14][54] = 8'hF4;
    assign wout[14][55] = 8'h02;
    assign wout[14][56] = 8'h10;
    assign wout[14][57] = 8'h1E;
    assign wout[14][58] = 8'h2C;
    assign wout[14][59] = 8'h3A;
    assign wout[14][60] = 8'h48;
    assign wout[14][61] = 8'h56;
    assign wout[14][62] = 8'h64;
    assign wout[14][63] = 8'h72;
    assign wout[15][0] = 8'h00;
    assign wout[15][1] = 8'h0F;
    assign wout[15][2] = 8'h1E;
    assign wout[15][3] = 8'h2D;
    assign wout[15][4] = 8'h3C;
    assign wout[15][5] = 8'h4B;
    assign wout[15][6] = 8'h5A;
    assign wout[15][7] = 8'h69;
    assign wout[15][8] = 8'h78;
    assign wout[15][9] = 8'h87;
    assign wout[15][10] = 8'h96;
    assign wout[15][11] = 8'hA5;
    assign wout[15][12] = 8'hB4;
    assign wout[15][13] = 8'hC3;
    assign wout[15][14] = 8'hD2;
    assign wout[15][15] = 8'hE1;
    assign wout[15][16] = 8'hF0;
    assign wout[15][17] = 8'hFF;
    assign wout[15][18] = 8'h0E;
    assign wout[15][19] = 8'h1D;
    assign wout[15][20] = 8'h2C;
    assign wout[15][21] = 8'h3B;
    assign wout[15][22] = 8'h4A;
    assign wout[15][23] = 8'h59;
    assign wout[15][24] = 8'h68;
    assign wout[15][25] = 8'h77;
    assign wout[15][26] = 8'h86;
    assign wout[15][27] = 8'h95;
    assign wout[15][28] = 8'hA4;
    assign wout[15][29] = 8'hB3;
    assign wout[15][30] = 8'hC2;
    assign wout[15][31] = 8'hD1;
    assign wout[15][32] = 8'hE0;
    assign wout[15][33] = 8'hEF;
    assign wout[15][34] = 8'hFE;
    assign wout[15][35] = 8'h0D;
    assign wout[15][36] = 8'h1C;
    assign wout[15][37] = 8'h2B;
    assign wout[15][38] = 8'h3A;
    assign wout[15][39] = 8'h49;
    assign wout[15][40] = 8'h58;
    assign wout[15][41] = 8'h67;
    assign wout[15][42] = 8'h76;
    assign wout[15][43] = 8'h85;
    assign wout[15][44] = 8'h94;
    assign wout[15][45] = 8'hA3;
    assign wout[15][46] = 8'hB2;
    assign wout[15][47] = 8'hC1;
    assign wout[15][48] = 8'hD0;
    assign wout[15][49] = 8'hDF;
    assign wout[15][50] = 8'hEE;
    assign wout[15][51] = 8'hFD;
    assign wout[15][52] = 8'h0C;
    assign wout[15][53] = 8'h1B;
    assign wout[15][54] = 8'h2A;
    assign wout[15][55] = 8'h39;
    assign wout[15][56] = 8'h48;
    assign wout[15][57] = 8'h57;
    assign wout[15][58] = 8'h66;
    assign wout[15][59] = 8'h75;
    assign wout[15][60] = 8'h84;
    assign wout[15][61] = 8'h93;
    assign wout[15][62] = 8'hA2;
    assign wout[15][63] = 8'hB1;
    assign wout[16][0] = 8'h00;
    assign wout[16][1] = 8'h10;
    assign wout[16][2] = 8'h20;
    assign wout[16][3] = 8'h30;
    assign wout[16][4] = 8'h40;
    assign wout[16][5] = 8'h50;
    assign wout[16][6] = 8'h60;
    assign wout[16][7] = 8'h70;
    assign wout[16][8] = 8'h80;
    assign wout[16][9] = 8'h90;
    assign wout[16][10] = 8'hA0;
    assign wout[16][11] = 8'hB0;
    assign wout[16][12] = 8'hC0;
    assign wout[16][13] = 8'hD0;
    assign wout[16][14] = 8'hE0;
    assign wout[16][15] = 8'hF0;
    assign wout[16][16] = 8'h00;
    assign wout[16][17] = 8'h10;
    assign wout[16][18] = 8'h20;
    assign wout[16][19] = 8'h30;
    assign wout[16][20] = 8'h40;
    assign wout[16][21] = 8'h50;
    assign wout[16][22] = 8'h60;
    assign wout[16][23] = 8'h70;
    assign wout[16][24] = 8'h80;
    assign wout[16][25] = 8'h90;
    assign wout[16][26] = 8'hA0;
    assign wout[16][27] = 8'hB0;
    assign wout[16][28] = 8'hC0;
    assign wout[16][29] = 8'hD0;
    assign wout[16][30] = 8'hE0;
    assign wout[16][31] = 8'hF0;
    assign wout[16][32] = 8'h00;
    assign wout[16][33] = 8'h10;
    assign wout[16][34] = 8'h20;
    assign wout[16][35] = 8'h30;
    assign wout[16][36] = 8'h40;
    assign wout[16][37] = 8'h50;
    assign wout[16][38] = 8'h60;
    assign wout[16][39] = 8'h70;
    assign wout[16][40] = 8'h80;
    assign wout[16][41] = 8'h90;
    assign wout[16][42] = 8'hA0;
    assign wout[16][43] = 8'hB0;
    assign wout[16][44] = 8'hC0;
    assign wout[16][45] = 8'hD0;
    assign wout[16][46] = 8'hE0;
    assign wout[16][47] = 8'hF0;
    assign wout[16][48] = 8'h00;
    assign wout[16][49] = 8'h10;
    assign wout[16][50] = 8'h20;
    assign wout[16][51] = 8'h30;
    assign wout[16][52] = 8'h40;
    assign wout[16][53] = 8'h50;
    assign wout[16][54] = 8'h60;
    assign wout[16][55] = 8'h70;
    assign wout[16][56] = 8'h80;
    assign wout[16][57] = 8'h90;
    assign wout[16][58] = 8'hA0;
    assign wout[16][59] = 8'hB0;
    assign wout[16][60] = 8'hC0;
    assign wout[16][61] = 8'hD0;
    assign wout[16][62] = 8'hE0;
    assign wout[16][63] = 8'hF0;
    assign wout[17][0] = 8'h00;
    assign wout[17][1] = 8'h11;
    assign wout[17][2] = 8'h22;
    assign wout[17][3] = 8'h33;
    assign wout[17][4] = 8'h44;
    assign wout[17][5] = 8'h55;
    assign wout[17][6] = 8'h66;
    assign wout[17][7] = 8'h77;
    assign wout[17][8] = 8'h88;
    assign wout[17][9] = 8'h99;
    assign wout[17][10] = 8'hAA;
    assign wout[17][11] = 8'hBB;
    assign wout[17][12] = 8'hCC;
    assign wout[17][13] = 8'hDD;
    assign wout[17][14] = 8'hEE;
    assign wout[17][15] = 8'hFF;
    assign wout[17][16] = 8'h10;
    assign wout[17][17] = 8'h21;
    assign wout[17][18] = 8'h32;
    assign wout[17][19] = 8'h43;
    assign wout[17][20] = 8'h54;
    assign wout[17][21] = 8'h65;
    assign wout[17][22] = 8'h76;
    assign wout[17][23] = 8'h87;
    assign wout[17][24] = 8'h98;
    assign wout[17][25] = 8'hA9;
    assign wout[17][26] = 8'hBA;
    assign wout[17][27] = 8'hCB;
    assign wout[17][28] = 8'hDC;
    assign wout[17][29] = 8'hED;
    assign wout[17][30] = 8'hFE;
    assign wout[17][31] = 8'h0F;
    assign wout[17][32] = 8'h20;
    assign wout[17][33] = 8'h31;
    assign wout[17][34] = 8'h42;
    assign wout[17][35] = 8'h53;
    assign wout[17][36] = 8'h64;
    assign wout[17][37] = 8'h75;
    assign wout[17][38] = 8'h86;
    assign wout[17][39] = 8'h97;
    assign wout[17][40] = 8'hA8;
    assign wout[17][41] = 8'hB9;
    assign wout[17][42] = 8'hCA;
    assign wout[17][43] = 8'hDB;
    assign wout[17][44] = 8'hEC;
    assign wout[17][45] = 8'hFD;
    assign wout[17][46] = 8'h0E;
    assign wout[17][47] = 8'h1F;
    assign wout[17][48] = 8'h30;
    assign wout[17][49] = 8'h41;
    assign wout[17][50] = 8'h52;
    assign wout[17][51] = 8'h63;
    assign wout[17][52] = 8'h74;
    assign wout[17][53] = 8'h85;
    assign wout[17][54] = 8'h96;
    assign wout[17][55] = 8'hA7;
    assign wout[17][56] = 8'hB8;
    assign wout[17][57] = 8'hC9;
    assign wout[17][58] = 8'hDA;
    assign wout[17][59] = 8'hEB;
    assign wout[17][60] = 8'hFC;
    assign wout[17][61] = 8'h0D;
    assign wout[17][62] = 8'h1E;
    assign wout[17][63] = 8'h2F;
    assign wout[18][0] = 8'h00;
    assign wout[18][1] = 8'h12;
    assign wout[18][2] = 8'h24;
    assign wout[18][3] = 8'h36;
    assign wout[18][4] = 8'h48;
    assign wout[18][5] = 8'h5A;
    assign wout[18][6] = 8'h6C;
    assign wout[18][7] = 8'h7E;
    assign wout[18][8] = 8'h90;
    assign wout[18][9] = 8'hA2;
    assign wout[18][10] = 8'hB4;
    assign wout[18][11] = 8'hC6;
    assign wout[18][12] = 8'hD8;
    assign wout[18][13] = 8'hEA;
    assign wout[18][14] = 8'hFC;
    assign wout[18][15] = 8'h0E;
    assign wout[18][16] = 8'h20;
    assign wout[18][17] = 8'h32;
    assign wout[18][18] = 8'h44;
    assign wout[18][19] = 8'h56;
    assign wout[18][20] = 8'h68;
    assign wout[18][21] = 8'h7A;
    assign wout[18][22] = 8'h8C;
    assign wout[18][23] = 8'h9E;
    assign wout[18][24] = 8'hB0;
    assign wout[18][25] = 8'hC2;
    assign wout[18][26] = 8'hD4;
    assign wout[18][27] = 8'hE6;
    assign wout[18][28] = 8'hF8;
    assign wout[18][29] = 8'h0A;
    assign wout[18][30] = 8'h1C;
    assign wout[18][31] = 8'h2E;
    assign wout[18][32] = 8'h40;
    assign wout[18][33] = 8'h52;
    assign wout[18][34] = 8'h64;
    assign wout[18][35] = 8'h76;
    assign wout[18][36] = 8'h88;
    assign wout[18][37] = 8'h9A;
    assign wout[18][38] = 8'hAC;
    assign wout[18][39] = 8'hBE;
    assign wout[18][40] = 8'hD0;
    assign wout[18][41] = 8'hE2;
    assign wout[18][42] = 8'hF4;
    assign wout[18][43] = 8'h06;
    assign wout[18][44] = 8'h18;
    assign wout[18][45] = 8'h2A;
    assign wout[18][46] = 8'h3C;
    assign wout[18][47] = 8'h4E;
    assign wout[18][48] = 8'h60;
    assign wout[18][49] = 8'h72;
    assign wout[18][50] = 8'h84;
    assign wout[18][51] = 8'h96;
    assign wout[18][52] = 8'hA8;
    assign wout[18][53] = 8'hBA;
    assign wout[18][54] = 8'hCC;
    assign wout[18][55] = 8'hDE;
    assign wout[18][56] = 8'hF0;
    assign wout[18][57] = 8'h02;
    assign wout[18][58] = 8'h14;
    assign wout[18][59] = 8'h26;
    assign wout[18][60] = 8'h38;
    assign wout[18][61] = 8'h4A;
    assign wout[18][62] = 8'h5C;
    assign wout[18][63] = 8'h6E;
    assign wout[19][0] = 8'h00;
    assign wout[19][1] = 8'h13;
    assign wout[19][2] = 8'h26;
    assign wout[19][3] = 8'h39;
    assign wout[19][4] = 8'h4C;
    assign wout[19][5] = 8'h5F;
    assign wout[19][6] = 8'h72;
    assign wout[19][7] = 8'h85;
    assign wout[19][8] = 8'h98;
    assign wout[19][9] = 8'hAB;
    assign wout[19][10] = 8'hBE;
    assign wout[19][11] = 8'hD1;
    assign wout[19][12] = 8'hE4;
    assign wout[19][13] = 8'hF7;
    assign wout[19][14] = 8'h0A;
    assign wout[19][15] = 8'h1D;
    assign wout[19][16] = 8'h30;
    assign wout[19][17] = 8'h43;
    assign wout[19][18] = 8'h56;
    assign wout[19][19] = 8'h69;
    assign wout[19][20] = 8'h7C;
    assign wout[19][21] = 8'h8F;
    assign wout[19][22] = 8'hA2;
    assign wout[19][23] = 8'hB5;
    assign wout[19][24] = 8'hC8;
    assign wout[19][25] = 8'hDB;
    assign wout[19][26] = 8'hEE;
    assign wout[19][27] = 8'h01;
    assign wout[19][28] = 8'h14;
    assign wout[19][29] = 8'h27;
    assign wout[19][30] = 8'h3A;
    assign wout[19][31] = 8'h4D;
    assign wout[19][32] = 8'h60;
    assign wout[19][33] = 8'h73;
    assign wout[19][34] = 8'h86;
    assign wout[19][35] = 8'h99;
    assign wout[19][36] = 8'hAC;
    assign wout[19][37] = 8'hBF;
    assign wout[19][38] = 8'hD2;
    assign wout[19][39] = 8'hE5;
    assign wout[19][40] = 8'hF8;
    assign wout[19][41] = 8'h0B;
    assign wout[19][42] = 8'h1E;
    assign wout[19][43] = 8'h31;
    assign wout[19][44] = 8'h44;
    assign wout[19][45] = 8'h57;
    assign wout[19][46] = 8'h6A;
    assign wout[19][47] = 8'h7D;
    assign wout[19][48] = 8'h90;
    assign wout[19][49] = 8'hA3;
    assign wout[19][50] = 8'hB6;
    assign wout[19][51] = 8'hC9;
    assign wout[19][52] = 8'hDC;
    assign wout[19][53] = 8'hEF;
    assign wout[19][54] = 8'h02;
    assign wout[19][55] = 8'h15;
    assign wout[19][56] = 8'h28;
    assign wout[19][57] = 8'h3B;
    assign wout[19][58] = 8'h4E;
    assign wout[19][59] = 8'h61;
    assign wout[19][60] = 8'h74;
    assign wout[19][61] = 8'h87;
    assign wout[19][62] = 8'h9A;
    assign wout[19][63] = 8'hAD;
    assign wout[20][0] = 8'h00;
    assign wout[20][1] = 8'h14;
    assign wout[20][2] = 8'h28;
    assign wout[20][3] = 8'h3C;
    assign wout[20][4] = 8'h50;
    assign wout[20][5] = 8'h64;
    assign wout[20][6] = 8'h78;
    assign wout[20][7] = 8'h8C;
    assign wout[20][8] = 8'hA0;
    assign wout[20][9] = 8'hB4;
    assign wout[20][10] = 8'hC8;
    assign wout[20][11] = 8'hDC;
    assign wout[20][12] = 8'hF0;
    assign wout[20][13] = 8'h04;
    assign wout[20][14] = 8'h18;
    assign wout[20][15] = 8'h2C;
    assign wout[20][16] = 8'h40;
    assign wout[20][17] = 8'h54;
    assign wout[20][18] = 8'h68;
    assign wout[20][19] = 8'h7C;
    assign wout[20][20] = 8'h90;
    assign wout[20][21] = 8'hA4;
    assign wout[20][22] = 8'hB8;
    assign wout[20][23] = 8'hCC;
    assign wout[20][24] = 8'hE0;
    assign wout[20][25] = 8'hF4;
    assign wout[20][26] = 8'h08;
    assign wout[20][27] = 8'h1C;
    assign wout[20][28] = 8'h30;
    assign wout[20][29] = 8'h44;
    assign wout[20][30] = 8'h58;
    assign wout[20][31] = 8'h6C;
    assign wout[20][32] = 8'h80;
    assign wout[20][33] = 8'h94;
    assign wout[20][34] = 8'hA8;
    assign wout[20][35] = 8'hBC;
    assign wout[20][36] = 8'hD0;
    assign wout[20][37] = 8'hE4;
    assign wout[20][38] = 8'hF8;
    assign wout[20][39] = 8'h0C;
    assign wout[20][40] = 8'h20;
    assign wout[20][41] = 8'h34;
    assign wout[20][42] = 8'h48;
    assign wout[20][43] = 8'h5C;
    assign wout[20][44] = 8'h70;
    assign wout[20][45] = 8'h84;
    assign wout[20][46] = 8'h98;
    assign wout[20][47] = 8'hAC;
    assign wout[20][48] = 8'hC0;
    assign wout[20][49] = 8'hD4;
    assign wout[20][50] = 8'hE8;
    assign wout[20][51] = 8'hFC;
    assign wout[20][52] = 8'h10;
    assign wout[20][53] = 8'h24;
    assign wout[20][54] = 8'h38;
    assign wout[20][55] = 8'h4C;
    assign wout[20][56] = 8'h60;
    assign wout[20][57] = 8'h74;
    assign wout[20][58] = 8'h88;
    assign wout[20][59] = 8'h9C;
    assign wout[20][60] = 8'hB0;
    assign wout[20][61] = 8'hC4;
    assign wout[20][62] = 8'hD8;
    assign wout[20][63] = 8'hEC;
    assign wout[21][0] = 8'h00;
    assign wout[21][1] = 8'h15;
    assign wout[21][2] = 8'h2A;
    assign wout[21][3] = 8'h3F;
    assign wout[21][4] = 8'h54;
    assign wout[21][5] = 8'h69;
    assign wout[21][6] = 8'h7E;
    assign wout[21][7] = 8'h93;
    assign wout[21][8] = 8'hA8;
    assign wout[21][9] = 8'hBD;
    assign wout[21][10] = 8'hD2;
    assign wout[21][11] = 8'hE7;
    assign wout[21][12] = 8'hFC;
    assign wout[21][13] = 8'h11;
    assign wout[21][14] = 8'h26;
    assign wout[21][15] = 8'h3B;
    assign wout[21][16] = 8'h50;
    assign wout[21][17] = 8'h65;
    assign wout[21][18] = 8'h7A;
    assign wout[21][19] = 8'h8F;
    assign wout[21][20] = 8'hA4;
    assign wout[21][21] = 8'hB9;
    assign wout[21][22] = 8'hCE;
    assign wout[21][23] = 8'hE3;
    assign wout[21][24] = 8'hF8;
    assign wout[21][25] = 8'h0D;
    assign wout[21][26] = 8'h22;
    assign wout[21][27] = 8'h37;
    assign wout[21][28] = 8'h4C;
    assign wout[21][29] = 8'h61;
    assign wout[21][30] = 8'h76;
    assign wout[21][31] = 8'h8B;
    assign wout[21][32] = 8'hA0;
    assign wout[21][33] = 8'hB5;
    assign wout[21][34] = 8'hCA;
    assign wout[21][35] = 8'hDF;
    assign wout[21][36] = 8'hF4;
    assign wout[21][37] = 8'h09;
    assign wout[21][38] = 8'h1E;
    assign wout[21][39] = 8'h33;
    assign wout[21][40] = 8'h48;
    assign wout[21][41] = 8'h5D;
    assign wout[21][42] = 8'h72;
    assign wout[21][43] = 8'h87;
    assign wout[21][44] = 8'h9C;
    assign wout[21][45] = 8'hB1;
    assign wout[21][46] = 8'hC6;
    assign wout[21][47] = 8'hDB;
    assign wout[21][48] = 8'hF0;
    assign wout[21][49] = 8'h05;
    assign wout[21][50] = 8'h1A;
    assign wout[21][51] = 8'h2F;
    assign wout[21][52] = 8'h44;
    assign wout[21][53] = 8'h59;
    assign wout[21][54] = 8'h6E;
    assign wout[21][55] = 8'h83;
    assign wout[21][56] = 8'h98;
    assign wout[21][57] = 8'hAD;
    assign wout[21][58] = 8'hC2;
    assign wout[21][59] = 8'hD7;
    assign wout[21][60] = 8'hEC;
    assign wout[21][61] = 8'h01;
    assign wout[21][62] = 8'h16;
    assign wout[21][63] = 8'h2B;
    assign wout[22][0] = 8'h00;
    assign wout[22][1] = 8'h16;
    assign wout[22][2] = 8'h2C;
    assign wout[22][3] = 8'h42;
    assign wout[22][4] = 8'h58;
    assign wout[22][5] = 8'h6E;
    assign wout[22][6] = 8'h84;
    assign wout[22][7] = 8'h9A;
    assign wout[22][8] = 8'hB0;
    assign wout[22][9] = 8'hC6;
    assign wout[22][10] = 8'hDC;
    assign wout[22][11] = 8'hF2;
    assign wout[22][12] = 8'h08;
    assign wout[22][13] = 8'h1E;
    assign wout[22][14] = 8'h34;
    assign wout[22][15] = 8'h4A;
    assign wout[22][16] = 8'h60;
    assign wout[22][17] = 8'h76;
    assign wout[22][18] = 8'h8C;
    assign wout[22][19] = 8'hA2;
    assign wout[22][20] = 8'hB8;
    assign wout[22][21] = 8'hCE;
    assign wout[22][22] = 8'hE4;
    assign wout[22][23] = 8'hFA;
    assign wout[22][24] = 8'h10;
    assign wout[22][25] = 8'h26;
    assign wout[22][26] = 8'h3C;
    assign wout[22][27] = 8'h52;
    assign wout[22][28] = 8'h68;
    assign wout[22][29] = 8'h7E;
    assign wout[22][30] = 8'h94;
    assign wout[22][31] = 8'hAA;
    assign wout[22][32] = 8'hC0;
    assign wout[22][33] = 8'hD6;
    assign wout[22][34] = 8'hEC;
    assign wout[22][35] = 8'h02;
    assign wout[22][36] = 8'h18;
    assign wout[22][37] = 8'h2E;
    assign wout[22][38] = 8'h44;
    assign wout[22][39] = 8'h5A;
    assign wout[22][40] = 8'h70;
    assign wout[22][41] = 8'h86;
    assign wout[22][42] = 8'h9C;
    assign wout[22][43] = 8'hB2;
    assign wout[22][44] = 8'hC8;
    assign wout[22][45] = 8'hDE;
    assign wout[22][46] = 8'hF4;
    assign wout[22][47] = 8'h0A;
    assign wout[22][48] = 8'h20;
    assign wout[22][49] = 8'h36;
    assign wout[22][50] = 8'h4C;
    assign wout[22][51] = 8'h62;
    assign wout[22][52] = 8'h78;
    assign wout[22][53] = 8'h8E;
    assign wout[22][54] = 8'hA4;
    assign wout[22][55] = 8'hBA;
    assign wout[22][56] = 8'hD0;
    assign wout[22][57] = 8'hE6;
    assign wout[22][58] = 8'hFC;
    assign wout[22][59] = 8'h12;
    assign wout[22][60] = 8'h28;
    assign wout[22][61] = 8'h3E;
    assign wout[22][62] = 8'h54;
    assign wout[22][63] = 8'h6A;
    assign wout[23][0] = 8'h00;
    assign wout[23][1] = 8'h17;
    assign wout[23][2] = 8'h2E;
    assign wout[23][3] = 8'h45;
    assign wout[23][4] = 8'h5C;
    assign wout[23][5] = 8'h73;
    assign wout[23][6] = 8'h8A;
    assign wout[23][7] = 8'hA1;
    assign wout[23][8] = 8'hB8;
    assign wout[23][9] = 8'hCF;
    assign wout[23][10] = 8'hE6;
    assign wout[23][11] = 8'hFD;
    assign wout[23][12] = 8'h14;
    assign wout[23][13] = 8'h2B;
    assign wout[23][14] = 8'h42;
    assign wout[23][15] = 8'h59;
    assign wout[23][16] = 8'h70;
    assign wout[23][17] = 8'h87;
    assign wout[23][18] = 8'h9E;
    assign wout[23][19] = 8'hB5;
    assign wout[23][20] = 8'hCC;
    assign wout[23][21] = 8'hE3;
    assign wout[23][22] = 8'hFA;
    assign wout[23][23] = 8'h11;
    assign wout[23][24] = 8'h28;
    assign wout[23][25] = 8'h3F;
    assign wout[23][26] = 8'h56;
    assign wout[23][27] = 8'h6D;
    assign wout[23][28] = 8'h84;
    assign wout[23][29] = 8'h9B;
    assign wout[23][30] = 8'hB2;
    assign wout[23][31] = 8'hC9;
    assign wout[23][32] = 8'hE0;
    assign wout[23][33] = 8'hF7;
    assign wout[23][34] = 8'h0E;
    assign wout[23][35] = 8'h25;
    assign wout[23][36] = 8'h3C;
    assign wout[23][37] = 8'h53;
    assign wout[23][38] = 8'h6A;
    assign wout[23][39] = 8'h81;
    assign wout[23][40] = 8'h98;
    assign wout[23][41] = 8'hAF;
    assign wout[23][42] = 8'hC6;
    assign wout[23][43] = 8'hDD;
    assign wout[23][44] = 8'hF4;
    assign wout[23][45] = 8'h0B;
    assign wout[23][46] = 8'h22;
    assign wout[23][47] = 8'h39;
    assign wout[23][48] = 8'h50;
    assign wout[23][49] = 8'h67;
    assign wout[23][50] = 8'h7E;
    assign wout[23][51] = 8'h95;
    assign wout[23][52] = 8'hAC;
    assign wout[23][53] = 8'hC3;
    assign wout[23][54] = 8'hDA;
    assign wout[23][55] = 8'hF1;
    assign wout[23][56] = 8'h08;
    assign wout[23][57] = 8'h1F;
    assign wout[23][58] = 8'h36;
    assign wout[23][59] = 8'h4D;
    assign wout[23][60] = 8'h64;
    assign wout[23][61] = 8'h7B;
    assign wout[23][62] = 8'h92;
    assign wout[23][63] = 8'hA9;
    assign wout[24][0] = 8'h00;
    assign wout[24][1] = 8'h18;
    assign wout[24][2] = 8'h30;
    assign wout[24][3] = 8'h48;
    assign wout[24][4] = 8'h60;
    assign wout[24][5] = 8'h78;
    assign wout[24][6] = 8'h90;
    assign wout[24][7] = 8'hA8;
    assign wout[24][8] = 8'hC0;
    assign wout[24][9] = 8'hD8;
    assign wout[24][10] = 8'hF0;
    assign wout[24][11] = 8'h08;
    assign wout[24][12] = 8'h20;
    assign wout[24][13] = 8'h38;
    assign wout[24][14] = 8'h50;
    assign wout[24][15] = 8'h68;
    assign wout[24][16] = 8'h80;
    assign wout[24][17] = 8'h98;
    assign wout[24][18] = 8'hB0;
    assign wout[24][19] = 8'hC8;
    assign wout[24][20] = 8'hE0;
    assign wout[24][21] = 8'hF8;
    assign wout[24][22] = 8'h10;
    assign wout[24][23] = 8'h28;
    assign wout[24][24] = 8'h40;
    assign wout[24][25] = 8'h58;
    assign wout[24][26] = 8'h70;
    assign wout[24][27] = 8'h88;
    assign wout[24][28] = 8'hA0;
    assign wout[24][29] = 8'hB8;
    assign wout[24][30] = 8'hD0;
    assign wout[24][31] = 8'hE8;
    assign wout[24][32] = 8'h00;
    assign wout[24][33] = 8'h18;
    assign wout[24][34] = 8'h30;
    assign wout[24][35] = 8'h48;
    assign wout[24][36] = 8'h60;
    assign wout[24][37] = 8'h78;
    assign wout[24][38] = 8'h90;
    assign wout[24][39] = 8'hA8;
    assign wout[24][40] = 8'hC0;
    assign wout[24][41] = 8'hD8;
    assign wout[24][42] = 8'hF0;
    assign wout[24][43] = 8'h08;
    assign wout[24][44] = 8'h20;
    assign wout[24][45] = 8'h38;
    assign wout[24][46] = 8'h50;
    assign wout[24][47] = 8'h68;
    assign wout[24][48] = 8'h80;
    assign wout[24][49] = 8'h98;
    assign wout[24][50] = 8'hB0;
    assign wout[24][51] = 8'hC8;
    assign wout[24][52] = 8'hE0;
    assign wout[24][53] = 8'hF8;
    assign wout[24][54] = 8'h10;
    assign wout[24][55] = 8'h28;
    assign wout[24][56] = 8'h40;
    assign wout[24][57] = 8'h58;
    assign wout[24][58] = 8'h70;
    assign wout[24][59] = 8'h88;
    assign wout[24][60] = 8'hA0;
    assign wout[24][61] = 8'hB8;
    assign wout[24][62] = 8'hD0;
    assign wout[24][63] = 8'hE8;
    assign wout[25][0] = 8'h00;
    assign wout[25][1] = 8'h19;
    assign wout[25][2] = 8'h32;
    assign wout[25][3] = 8'h4B;
    assign wout[25][4] = 8'h64;
    assign wout[25][5] = 8'h7D;
    assign wout[25][6] = 8'h96;
    assign wout[25][7] = 8'hAF;
    assign wout[25][8] = 8'hC8;
    assign wout[25][9] = 8'hE1;
    assign wout[25][10] = 8'hFA;
    assign wout[25][11] = 8'h13;
    assign wout[25][12] = 8'h2C;
    assign wout[25][13] = 8'h45;
    assign wout[25][14] = 8'h5E;
    assign wout[25][15] = 8'h77;
    assign wout[25][16] = 8'h90;
    assign wout[25][17] = 8'hA9;
    assign wout[25][18] = 8'hC2;
    assign wout[25][19] = 8'hDB;
    assign wout[25][20] = 8'hF4;
    assign wout[25][21] = 8'h0D;
    assign wout[25][22] = 8'h26;
    assign wout[25][23] = 8'h3F;
    assign wout[25][24] = 8'h58;
    assign wout[25][25] = 8'h71;
    assign wout[25][26] = 8'h8A;
    assign wout[25][27] = 8'hA3;
    assign wout[25][28] = 8'hBC;
    assign wout[25][29] = 8'hD5;
    assign wout[25][30] = 8'hEE;
    assign wout[25][31] = 8'h07;
    assign wout[25][32] = 8'h20;
    assign wout[25][33] = 8'h39;
    assign wout[25][34] = 8'h52;
    assign wout[25][35] = 8'h6B;
    assign wout[25][36] = 8'h84;
    assign wout[25][37] = 8'h9D;
    assign wout[25][38] = 8'hB6;
    assign wout[25][39] = 8'hCF;
    assign wout[25][40] = 8'hE8;
    assign wout[25][41] = 8'h01;
    assign wout[25][42] = 8'h1A;
    assign wout[25][43] = 8'h33;
    assign wout[25][44] = 8'h4C;
    assign wout[25][45] = 8'h65;
    assign wout[25][46] = 8'h7E;
    assign wout[25][47] = 8'h97;
    assign wout[25][48] = 8'hB0;
    assign wout[25][49] = 8'hC9;
    assign wout[25][50] = 8'hE2;
    assign wout[25][51] = 8'hFB;
    assign wout[25][52] = 8'h14;
    assign wout[25][53] = 8'h2D;
    assign wout[25][54] = 8'h46;
    assign wout[25][55] = 8'h5F;
    assign wout[25][56] = 8'h78;
    assign wout[25][57] = 8'h91;
    assign wout[25][58] = 8'hAA;
    assign wout[25][59] = 8'hC3;
    assign wout[25][60] = 8'hDC;
    assign wout[25][61] = 8'hF5;
    assign wout[25][62] = 8'h0E;
    assign wout[25][63] = 8'h27;
    assign wout[26][0] = 8'h00;
    assign wout[26][1] = 8'h1A;
    assign wout[26][2] = 8'h34;
    assign wout[26][3] = 8'h4E;
    assign wout[26][4] = 8'h68;
    assign wout[26][5] = 8'h82;
    assign wout[26][6] = 8'h9C;
    assign wout[26][7] = 8'hB6;
    assign wout[26][8] = 8'hD0;
    assign wout[26][9] = 8'hEA;
    assign wout[26][10] = 8'h04;
    assign wout[26][11] = 8'h1E;
    assign wout[26][12] = 8'h38;
    assign wout[26][13] = 8'h52;
    assign wout[26][14] = 8'h6C;
    assign wout[26][15] = 8'h86;
    assign wout[26][16] = 8'hA0;
    assign wout[26][17] = 8'hBA;
    assign wout[26][18] = 8'hD4;
    assign wout[26][19] = 8'hEE;
    assign wout[26][20] = 8'h08;
    assign wout[26][21] = 8'h22;
    assign wout[26][22] = 8'h3C;
    assign wout[26][23] = 8'h56;
    assign wout[26][24] = 8'h70;
    assign wout[26][25] = 8'h8A;
    assign wout[26][26] = 8'hA4;
    assign wout[26][27] = 8'hBE;
    assign wout[26][28] = 8'hD8;
    assign wout[26][29] = 8'hF2;
    assign wout[26][30] = 8'h0C;
    assign wout[26][31] = 8'h26;
    assign wout[26][32] = 8'h40;
    assign wout[26][33] = 8'h5A;
    assign wout[26][34] = 8'h74;
    assign wout[26][35] = 8'h8E;
    assign wout[26][36] = 8'hA8;
    assign wout[26][37] = 8'hC2;
    assign wout[26][38] = 8'hDC;
    assign wout[26][39] = 8'hF6;
    assign wout[26][40] = 8'h10;
    assign wout[26][41] = 8'h2A;
    assign wout[26][42] = 8'h44;
    assign wout[26][43] = 8'h5E;
    assign wout[26][44] = 8'h78;
    assign wout[26][45] = 8'h92;
    assign wout[26][46] = 8'hAC;
    assign wout[26][47] = 8'hC6;
    assign wout[26][48] = 8'hE0;
    assign wout[26][49] = 8'hFA;
    assign wout[26][50] = 8'h14;
    assign wout[26][51] = 8'h2E;
    assign wout[26][52] = 8'h48;
    assign wout[26][53] = 8'h62;
    assign wout[26][54] = 8'h7C;
    assign wout[26][55] = 8'h96;
    assign wout[26][56] = 8'hB0;
    assign wout[26][57] = 8'hCA;
    assign wout[26][58] = 8'hE4;
    assign wout[26][59] = 8'hFE;
    assign wout[26][60] = 8'h18;
    assign wout[26][61] = 8'h32;
    assign wout[26][62] = 8'h4C;
    assign wout[26][63] = 8'h66;
    assign wout[27][0] = 8'h00;
    assign wout[27][1] = 8'h1B;
    assign wout[27][2] = 8'h36;
    assign wout[27][3] = 8'h51;
    assign wout[27][4] = 8'h6C;
    assign wout[27][5] = 8'h87;
    assign wout[27][6] = 8'hA2;
    assign wout[27][7] = 8'hBD;
    assign wout[27][8] = 8'hD8;
    assign wout[27][9] = 8'hF3;
    assign wout[27][10] = 8'h0E;
    assign wout[27][11] = 8'h29;
    assign wout[27][12] = 8'h44;
    assign wout[27][13] = 8'h5F;
    assign wout[27][14] = 8'h7A;
    assign wout[27][15] = 8'h95;
    assign wout[27][16] = 8'hB0;
    assign wout[27][17] = 8'hCB;
    assign wout[27][18] = 8'hE6;
    assign wout[27][19] = 8'h01;
    assign wout[27][20] = 8'h1C;
    assign wout[27][21] = 8'h37;
    assign wout[27][22] = 8'h52;
    assign wout[27][23] = 8'h6D;
    assign wout[27][24] = 8'h88;
    assign wout[27][25] = 8'hA3;
    assign wout[27][26] = 8'hBE;
    assign wout[27][27] = 8'hD9;
    assign wout[27][28] = 8'hF4;
    assign wout[27][29] = 8'h0F;
    assign wout[27][30] = 8'h2A;
    assign wout[27][31] = 8'h45;
    assign wout[27][32] = 8'h60;
    assign wout[27][33] = 8'h7B;
    assign wout[27][34] = 8'h96;
    assign wout[27][35] = 8'hB1;
    assign wout[27][36] = 8'hCC;
    assign wout[27][37] = 8'hE7;
    assign wout[27][38] = 8'h02;
    assign wout[27][39] = 8'h1D;
    assign wout[27][40] = 8'h38;
    assign wout[27][41] = 8'h53;
    assign wout[27][42] = 8'h6E;
    assign wout[27][43] = 8'h89;
    assign wout[27][44] = 8'hA4;
    assign wout[27][45] = 8'hBF;
    assign wout[27][46] = 8'hDA;
    assign wout[27][47] = 8'hF5;
    assign wout[27][48] = 8'h10;
    assign wout[27][49] = 8'h2B;
    assign wout[27][50] = 8'h46;
    assign wout[27][51] = 8'h61;
    assign wout[27][52] = 8'h7C;
    assign wout[27][53] = 8'h97;
    assign wout[27][54] = 8'hB2;
    assign wout[27][55] = 8'hCD;
    assign wout[27][56] = 8'hE8;
    assign wout[27][57] = 8'h03;
    assign wout[27][58] = 8'h1E;
    assign wout[27][59] = 8'h39;
    assign wout[27][60] = 8'h54;
    assign wout[27][61] = 8'h6F;
    assign wout[27][62] = 8'h8A;
    assign wout[27][63] = 8'hA5;
    assign wout[28][0] = 8'h00;
    assign wout[28][1] = 8'h1C;
    assign wout[28][2] = 8'h38;
    assign wout[28][3] = 8'h54;
    assign wout[28][4] = 8'h70;
    assign wout[28][5] = 8'h8C;
    assign wout[28][6] = 8'hA8;
    assign wout[28][7] = 8'hC4;
    assign wout[28][8] = 8'hE0;
    assign wout[28][9] = 8'hFC;
    assign wout[28][10] = 8'h18;
    assign wout[28][11] = 8'h34;
    assign wout[28][12] = 8'h50;
    assign wout[28][13] = 8'h6C;
    assign wout[28][14] = 8'h88;
    assign wout[28][15] = 8'hA4;
    assign wout[28][16] = 8'hC0;
    assign wout[28][17] = 8'hDC;
    assign wout[28][18] = 8'hF8;
    assign wout[28][19] = 8'h14;
    assign wout[28][20] = 8'h30;
    assign wout[28][21] = 8'h4C;
    assign wout[28][22] = 8'h68;
    assign wout[28][23] = 8'h84;
    assign wout[28][24] = 8'hA0;
    assign wout[28][25] = 8'hBC;
    assign wout[28][26] = 8'hD8;
    assign wout[28][27] = 8'hF4;
    assign wout[28][28] = 8'h10;
    assign wout[28][29] = 8'h2C;
    assign wout[28][30] = 8'h48;
    assign wout[28][31] = 8'h64;
    assign wout[28][32] = 8'h80;
    assign wout[28][33] = 8'h9C;
    assign wout[28][34] = 8'hB8;
    assign wout[28][35] = 8'hD4;
    assign wout[28][36] = 8'hF0;
    assign wout[28][37] = 8'h0C;
    assign wout[28][38] = 8'h28;
    assign wout[28][39] = 8'h44;
    assign wout[28][40] = 8'h60;
    assign wout[28][41] = 8'h7C;
    assign wout[28][42] = 8'h98;
    assign wout[28][43] = 8'hB4;
    assign wout[28][44] = 8'hD0;
    assign wout[28][45] = 8'hEC;
    assign wout[28][46] = 8'h08;
    assign wout[28][47] = 8'h24;
    assign wout[28][48] = 8'h40;
    assign wout[28][49] = 8'h5C;
    assign wout[28][50] = 8'h78;
    assign wout[28][51] = 8'h94;
    assign wout[28][52] = 8'hB0;
    assign wout[28][53] = 8'hCC;
    assign wout[28][54] = 8'hE8;
    assign wout[28][55] = 8'h04;
    assign wout[28][56] = 8'h20;
    assign wout[28][57] = 8'h3C;
    assign wout[28][58] = 8'h58;
    assign wout[28][59] = 8'h74;
    assign wout[28][60] = 8'h90;
    assign wout[28][61] = 8'hAC;
    assign wout[28][62] = 8'hC8;
    assign wout[28][63] = 8'hE4;
    assign wout[29][0] = 8'h00;
    assign wout[29][1] = 8'h1D;
    assign wout[29][2] = 8'h3A;
    assign wout[29][3] = 8'h57;
    assign wout[29][4] = 8'h74;
    assign wout[29][5] = 8'h91;
    assign wout[29][6] = 8'hAE;
    assign wout[29][7] = 8'hCB;
    assign wout[29][8] = 8'hE8;
    assign wout[29][9] = 8'h05;
    assign wout[29][10] = 8'h22;
    assign wout[29][11] = 8'h3F;
    assign wout[29][12] = 8'h5C;
    assign wout[29][13] = 8'h79;
    assign wout[29][14] = 8'h96;
    assign wout[29][15] = 8'hB3;
    assign wout[29][16] = 8'hD0;
    assign wout[29][17] = 8'hED;
    assign wout[29][18] = 8'h0A;
    assign wout[29][19] = 8'h27;
    assign wout[29][20] = 8'h44;
    assign wout[29][21] = 8'h61;
    assign wout[29][22] = 8'h7E;
    assign wout[29][23] = 8'h9B;
    assign wout[29][24] = 8'hB8;
    assign wout[29][25] = 8'hD5;
    assign wout[29][26] = 8'hF2;
    assign wout[29][27] = 8'h0F;
    assign wout[29][28] = 8'h2C;
    assign wout[29][29] = 8'h49;
    assign wout[29][30] = 8'h66;
    assign wout[29][31] = 8'h83;
    assign wout[29][32] = 8'hA0;
    assign wout[29][33] = 8'hBD;
    assign wout[29][34] = 8'hDA;
    assign wout[29][35] = 8'hF7;
    assign wout[29][36] = 8'h14;
    assign wout[29][37] = 8'h31;
    assign wout[29][38] = 8'h4E;
    assign wout[29][39] = 8'h6B;
    assign wout[29][40] = 8'h88;
    assign wout[29][41] = 8'hA5;
    assign wout[29][42] = 8'hC2;
    assign wout[29][43] = 8'hDF;
    assign wout[29][44] = 8'hFC;
    assign wout[29][45] = 8'h19;
    assign wout[29][46] = 8'h36;
    assign wout[29][47] = 8'h53;
    assign wout[29][48] = 8'h70;
    assign wout[29][49] = 8'h8D;
    assign wout[29][50] = 8'hAA;
    assign wout[29][51] = 8'hC7;
    assign wout[29][52] = 8'hE4;
    assign wout[29][53] = 8'h01;
    assign wout[29][54] = 8'h1E;
    assign wout[29][55] = 8'h3B;
    assign wout[29][56] = 8'h58;
    assign wout[29][57] = 8'h75;
    assign wout[29][58] = 8'h92;
    assign wout[29][59] = 8'hAF;
    assign wout[29][60] = 8'hCC;
    assign wout[29][61] = 8'hE9;
    assign wout[29][62] = 8'h06;
    assign wout[29][63] = 8'h23;
    assign wout[30][0] = 8'h00;
    assign wout[30][1] = 8'h1E;
    assign wout[30][2] = 8'h3C;
    assign wout[30][3] = 8'h5A;
    assign wout[30][4] = 8'h78;
    assign wout[30][5] = 8'h96;
    assign wout[30][6] = 8'hB4;
    assign wout[30][7] = 8'hD2;
    assign wout[30][8] = 8'hF0;
    assign wout[30][9] = 8'h0E;
    assign wout[30][10] = 8'h2C;
    assign wout[30][11] = 8'h4A;
    assign wout[30][12] = 8'h68;
    assign wout[30][13] = 8'h86;
    assign wout[30][14] = 8'hA4;
    assign wout[30][15] = 8'hC2;
    assign wout[30][16] = 8'hE0;
    assign wout[30][17] = 8'hFE;
    assign wout[30][18] = 8'h1C;
    assign wout[30][19] = 8'h3A;
    assign wout[30][20] = 8'h58;
    assign wout[30][21] = 8'h76;
    assign wout[30][22] = 8'h94;
    assign wout[30][23] = 8'hB2;
    assign wout[30][24] = 8'hD0;
    assign wout[30][25] = 8'hEE;
    assign wout[30][26] = 8'h0C;
    assign wout[30][27] = 8'h2A;
    assign wout[30][28] = 8'h48;
    assign wout[30][29] = 8'h66;
    assign wout[30][30] = 8'h84;
    assign wout[30][31] = 8'hA2;
    assign wout[30][32] = 8'hC0;
    assign wout[30][33] = 8'hDE;
    assign wout[30][34] = 8'hFC;
    assign wout[30][35] = 8'h1A;
    assign wout[30][36] = 8'h38;
    assign wout[30][37] = 8'h56;
    assign wout[30][38] = 8'h74;
    assign wout[30][39] = 8'h92;
    assign wout[30][40] = 8'hB0;
    assign wout[30][41] = 8'hCE;
    assign wout[30][42] = 8'hEC;
    assign wout[30][43] = 8'h0A;
    assign wout[30][44] = 8'h28;
    assign wout[30][45] = 8'h46;
    assign wout[30][46] = 8'h64;
    assign wout[30][47] = 8'h82;
    assign wout[30][48] = 8'hA0;
    assign wout[30][49] = 8'hBE;
    assign wout[30][50] = 8'hDC;
    assign wout[30][51] = 8'hFA;
    assign wout[30][52] = 8'h18;
    assign wout[30][53] = 8'h36;
    assign wout[30][54] = 8'h54;
    assign wout[30][55] = 8'h72;
    assign wout[30][56] = 8'h90;
    assign wout[30][57] = 8'hAE;
    assign wout[30][58] = 8'hCC;
    assign wout[30][59] = 8'hEA;
    assign wout[30][60] = 8'h08;
    assign wout[30][61] = 8'h26;
    assign wout[30][62] = 8'h44;
    assign wout[30][63] = 8'h62;
    assign wout[31][0] = 8'h00;
    assign wout[31][1] = 8'h1F;
    assign wout[31][2] = 8'h3E;
    assign wout[31][3] = 8'h5D;
    assign wout[31][4] = 8'h7C;
    assign wout[31][5] = 8'h9B;
    assign wout[31][6] = 8'hBA;
    assign wout[31][7] = 8'hD9;
    assign wout[31][8] = 8'hF8;
    assign wout[31][9] = 8'h17;
    assign wout[31][10] = 8'h36;
    assign wout[31][11] = 8'h55;
    assign wout[31][12] = 8'h74;
    assign wout[31][13] = 8'h93;
    assign wout[31][14] = 8'hB2;
    assign wout[31][15] = 8'hD1;
    assign wout[31][16] = 8'hF0;
    assign wout[31][17] = 8'h0F;
    assign wout[31][18] = 8'h2E;
    assign wout[31][19] = 8'h4D;
    assign wout[31][20] = 8'h6C;
    assign wout[31][21] = 8'h8B;
    assign wout[31][22] = 8'hAA;
    assign wout[31][23] = 8'hC9;
    assign wout[31][24] = 8'hE8;
    assign wout[31][25] = 8'h07;
    assign wout[31][26] = 8'h26;
    assign wout[31][27] = 8'h45;
    assign wout[31][28] = 8'h64;
    assign wout[31][29] = 8'h83;
    assign wout[31][30] = 8'hA2;
    assign wout[31][31] = 8'hC1;
    assign wout[31][32] = 8'hE0;
    assign wout[31][33] = 8'hFF;
    assign wout[31][34] = 8'h1E;
    assign wout[31][35] = 8'h3D;
    assign wout[31][36] = 8'h5C;
    assign wout[31][37] = 8'h7B;
    assign wout[31][38] = 8'h9A;
    assign wout[31][39] = 8'hB9;
    assign wout[31][40] = 8'hD8;
    assign wout[31][41] = 8'hF7;
    assign wout[31][42] = 8'h16;
    assign wout[31][43] = 8'h35;
    assign wout[31][44] = 8'h54;
    assign wout[31][45] = 8'h73;
    assign wout[31][46] = 8'h92;
    assign wout[31][47] = 8'hB1;
    assign wout[31][48] = 8'hD0;
    assign wout[31][49] = 8'hEF;
    assign wout[31][50] = 8'h0E;
    assign wout[31][51] = 8'h2D;
    assign wout[31][52] = 8'h4C;
    assign wout[31][53] = 8'h6B;
    assign wout[31][54] = 8'h8A;
    assign wout[31][55] = 8'hA9;
    assign wout[31][56] = 8'hC8;
    assign wout[31][57] = 8'hE7;
    assign wout[31][58] = 8'h06;
    assign wout[31][59] = 8'h25;
    assign wout[31][60] = 8'h44;
    assign wout[31][61] = 8'h63;
    assign wout[31][62] = 8'h82;
    assign wout[31][63] = 8'hA1;
    assign wout[32][0] = 8'h00;
    assign wout[32][1] = 8'h20;
    assign wout[32][2] = 8'h40;
    assign wout[32][3] = 8'h60;
    assign wout[32][4] = 8'h80;
    assign wout[32][5] = 8'hA0;
    assign wout[32][6] = 8'hC0;
    assign wout[32][7] = 8'hE0;
    assign wout[32][8] = 8'h00;
    assign wout[32][9] = 8'h20;
    assign wout[32][10] = 8'h40;
    assign wout[32][11] = 8'h60;
    assign wout[32][12] = 8'h80;
    assign wout[32][13] = 8'hA0;
    assign wout[32][14] = 8'hC0;
    assign wout[32][15] = 8'hE0;
    assign wout[32][16] = 8'h00;
    assign wout[32][17] = 8'h20;
    assign wout[32][18] = 8'h40;
    assign wout[32][19] = 8'h60;
    assign wout[32][20] = 8'h80;
    assign wout[32][21] = 8'hA0;
    assign wout[32][22] = 8'hC0;
    assign wout[32][23] = 8'hE0;
    assign wout[32][24] = 8'h00;
    assign wout[32][25] = 8'h20;
    assign wout[32][26] = 8'h40;
    assign wout[32][27] = 8'h60;
    assign wout[32][28] = 8'h80;
    assign wout[32][29] = 8'hA0;
    assign wout[32][30] = 8'hC0;
    assign wout[32][31] = 8'hE0;
    assign wout[32][32] = 8'h00;
    assign wout[32][33] = 8'h20;
    assign wout[32][34] = 8'h40;
    assign wout[32][35] = 8'h60;
    assign wout[32][36] = 8'h80;
    assign wout[32][37] = 8'hA0;
    assign wout[32][38] = 8'hC0;
    assign wout[32][39] = 8'hE0;
    assign wout[32][40] = 8'h00;
    assign wout[32][41] = 8'h20;
    assign wout[32][42] = 8'h40;
    assign wout[32][43] = 8'h60;
    assign wout[32][44] = 8'h80;
    assign wout[32][45] = 8'hA0;
    assign wout[32][46] = 8'hC0;
    assign wout[32][47] = 8'hE0;
    assign wout[32][48] = 8'h00;
    assign wout[32][49] = 8'h20;
    assign wout[32][50] = 8'h40;
    assign wout[32][51] = 8'h60;
    assign wout[32][52] = 8'h80;
    assign wout[32][53] = 8'hA0;
    assign wout[32][54] = 8'hC0;
    assign wout[32][55] = 8'hE0;
    assign wout[32][56] = 8'h00;
    assign wout[32][57] = 8'h20;
    assign wout[32][58] = 8'h40;
    assign wout[32][59] = 8'h60;
    assign wout[32][60] = 8'h80;
    assign wout[32][61] = 8'hA0;
    assign wout[32][62] = 8'hC0;
    assign wout[32][63] = 8'hE0;
    assign wout[33][0] = 8'h00;
    assign wout[33][1] = 8'h21;
    assign wout[33][2] = 8'h42;
    assign wout[33][3] = 8'h63;
    assign wout[33][4] = 8'h84;
    assign wout[33][5] = 8'hA5;
    assign wout[33][6] = 8'hC6;
    assign wout[33][7] = 8'hE7;
    assign wout[33][8] = 8'h08;
    assign wout[33][9] = 8'h29;
    assign wout[33][10] = 8'h4A;
    assign wout[33][11] = 8'h6B;
    assign wout[33][12] = 8'h8C;
    assign wout[33][13] = 8'hAD;
    assign wout[33][14] = 8'hCE;
    assign wout[33][15] = 8'hEF;
    assign wout[33][16] = 8'h10;
    assign wout[33][17] = 8'h31;
    assign wout[33][18] = 8'h52;
    assign wout[33][19] = 8'h73;
    assign wout[33][20] = 8'h94;
    assign wout[33][21] = 8'hB5;
    assign wout[33][22] = 8'hD6;
    assign wout[33][23] = 8'hF7;
    assign wout[33][24] = 8'h18;
    assign wout[33][25] = 8'h39;
    assign wout[33][26] = 8'h5A;
    assign wout[33][27] = 8'h7B;
    assign wout[33][28] = 8'h9C;
    assign wout[33][29] = 8'hBD;
    assign wout[33][30] = 8'hDE;
    assign wout[33][31] = 8'hFF;
    assign wout[33][32] = 8'h20;
    assign wout[33][33] = 8'h41;
    assign wout[33][34] = 8'h62;
    assign wout[33][35] = 8'h83;
    assign wout[33][36] = 8'hA4;
    assign wout[33][37] = 8'hC5;
    assign wout[33][38] = 8'hE6;
    assign wout[33][39] = 8'h07;
    assign wout[33][40] = 8'h28;
    assign wout[33][41] = 8'h49;
    assign wout[33][42] = 8'h6A;
    assign wout[33][43] = 8'h8B;
    assign wout[33][44] = 8'hAC;
    assign wout[33][45] = 8'hCD;
    assign wout[33][46] = 8'hEE;
    assign wout[33][47] = 8'h0F;
    assign wout[33][48] = 8'h30;
    assign wout[33][49] = 8'h51;
    assign wout[33][50] = 8'h72;
    assign wout[33][51] = 8'h93;
    assign wout[33][52] = 8'hB4;
    assign wout[33][53] = 8'hD5;
    assign wout[33][54] = 8'hF6;
    assign wout[33][55] = 8'h17;
    assign wout[33][56] = 8'h38;
    assign wout[33][57] = 8'h59;
    assign wout[33][58] = 8'h7A;
    assign wout[33][59] = 8'h9B;
    assign wout[33][60] = 8'hBC;
    assign wout[33][61] = 8'hDD;
    assign wout[33][62] = 8'hFE;
    assign wout[33][63] = 8'h1F;
    assign wout[34][0] = 8'h00;
    assign wout[34][1] = 8'h22;
    assign wout[34][2] = 8'h44;
    assign wout[34][3] = 8'h66;
    assign wout[34][4] = 8'h88;
    assign wout[34][5] = 8'hAA;
    assign wout[34][6] = 8'hCC;
    assign wout[34][7] = 8'hEE;
    assign wout[34][8] = 8'h10;
    assign wout[34][9] = 8'h32;
    assign wout[34][10] = 8'h54;
    assign wout[34][11] = 8'h76;
    assign wout[34][12] = 8'h98;
    assign wout[34][13] = 8'hBA;
    assign wout[34][14] = 8'hDC;
    assign wout[34][15] = 8'hFE;
    assign wout[34][16] = 8'h20;
    assign wout[34][17] = 8'h42;
    assign wout[34][18] = 8'h64;
    assign wout[34][19] = 8'h86;
    assign wout[34][20] = 8'hA8;
    assign wout[34][21] = 8'hCA;
    assign wout[34][22] = 8'hEC;
    assign wout[34][23] = 8'h0E;
    assign wout[34][24] = 8'h30;
    assign wout[34][25] = 8'h52;
    assign wout[34][26] = 8'h74;
    assign wout[34][27] = 8'h96;
    assign wout[34][28] = 8'hB8;
    assign wout[34][29] = 8'hDA;
    assign wout[34][30] = 8'hFC;
    assign wout[34][31] = 8'h1E;
    assign wout[34][32] = 8'h40;
    assign wout[34][33] = 8'h62;
    assign wout[34][34] = 8'h84;
    assign wout[34][35] = 8'hA6;
    assign wout[34][36] = 8'hC8;
    assign wout[34][37] = 8'hEA;
    assign wout[34][38] = 8'h0C;
    assign wout[34][39] = 8'h2E;
    assign wout[34][40] = 8'h50;
    assign wout[34][41] = 8'h72;
    assign wout[34][42] = 8'h94;
    assign wout[34][43] = 8'hB6;
    assign wout[34][44] = 8'hD8;
    assign wout[34][45] = 8'hFA;
    assign wout[34][46] = 8'h1C;
    assign wout[34][47] = 8'h3E;
    assign wout[34][48] = 8'h60;
    assign wout[34][49] = 8'h82;
    assign wout[34][50] = 8'hA4;
    assign wout[34][51] = 8'hC6;
    assign wout[34][52] = 8'hE8;
    assign wout[34][53] = 8'h0A;
    assign wout[34][54] = 8'h2C;
    assign wout[34][55] = 8'h4E;
    assign wout[34][56] = 8'h70;
    assign wout[34][57] = 8'h92;
    assign wout[34][58] = 8'hB4;
    assign wout[34][59] = 8'hD6;
    assign wout[34][60] = 8'hF8;
    assign wout[34][61] = 8'h1A;
    assign wout[34][62] = 8'h3C;
    assign wout[34][63] = 8'h5E;
    assign wout[35][0] = 8'h00;
    assign wout[35][1] = 8'h23;
    assign wout[35][2] = 8'h46;
    assign wout[35][3] = 8'h69;
    assign wout[35][4] = 8'h8C;
    assign wout[35][5] = 8'hAF;
    assign wout[35][6] = 8'hD2;
    assign wout[35][7] = 8'hF5;
    assign wout[35][8] = 8'h18;
    assign wout[35][9] = 8'h3B;
    assign wout[35][10] = 8'h5E;
    assign wout[35][11] = 8'h81;
    assign wout[35][12] = 8'hA4;
    assign wout[35][13] = 8'hC7;
    assign wout[35][14] = 8'hEA;
    assign wout[35][15] = 8'h0D;
    assign wout[35][16] = 8'h30;
    assign wout[35][17] = 8'h53;
    assign wout[35][18] = 8'h76;
    assign wout[35][19] = 8'h99;
    assign wout[35][20] = 8'hBC;
    assign wout[35][21] = 8'hDF;
    assign wout[35][22] = 8'h02;
    assign wout[35][23] = 8'h25;
    assign wout[35][24] = 8'h48;
    assign wout[35][25] = 8'h6B;
    assign wout[35][26] = 8'h8E;
    assign wout[35][27] = 8'hB1;
    assign wout[35][28] = 8'hD4;
    assign wout[35][29] = 8'hF7;
    assign wout[35][30] = 8'h1A;
    assign wout[35][31] = 8'h3D;
    assign wout[35][32] = 8'h60;
    assign wout[35][33] = 8'h83;
    assign wout[35][34] = 8'hA6;
    assign wout[35][35] = 8'hC9;
    assign wout[35][36] = 8'hEC;
    assign wout[35][37] = 8'h0F;
    assign wout[35][38] = 8'h32;
    assign wout[35][39] = 8'h55;
    assign wout[35][40] = 8'h78;
    assign wout[35][41] = 8'h9B;
    assign wout[35][42] = 8'hBE;
    assign wout[35][43] = 8'hE1;
    assign wout[35][44] = 8'h04;
    assign wout[35][45] = 8'h27;
    assign wout[35][46] = 8'h4A;
    assign wout[35][47] = 8'h6D;
    assign wout[35][48] = 8'h90;
    assign wout[35][49] = 8'hB3;
    assign wout[35][50] = 8'hD6;
    assign wout[35][51] = 8'hF9;
    assign wout[35][52] = 8'h1C;
    assign wout[35][53] = 8'h3F;
    assign wout[35][54] = 8'h62;
    assign wout[35][55] = 8'h85;
    assign wout[35][56] = 8'hA8;
    assign wout[35][57] = 8'hCB;
    assign wout[35][58] = 8'hEE;
    assign wout[35][59] = 8'h11;
    assign wout[35][60] = 8'h34;
    assign wout[35][61] = 8'h57;
    assign wout[35][62] = 8'h7A;
    assign wout[35][63] = 8'h9D;
    assign wout[36][0] = 8'h00;
    assign wout[36][1] = 8'h24;
    assign wout[36][2] = 8'h48;
    assign wout[36][3] = 8'h6C;
    assign wout[36][4] = 8'h90;
    assign wout[36][5] = 8'hB4;
    assign wout[36][6] = 8'hD8;
    assign wout[36][7] = 8'hFC;
    assign wout[36][8] = 8'h20;
    assign wout[36][9] = 8'h44;
    assign wout[36][10] = 8'h68;
    assign wout[36][11] = 8'h8C;
    assign wout[36][12] = 8'hB0;
    assign wout[36][13] = 8'hD4;
    assign wout[36][14] = 8'hF8;
    assign wout[36][15] = 8'h1C;
    assign wout[36][16] = 8'h40;
    assign wout[36][17] = 8'h64;
    assign wout[36][18] = 8'h88;
    assign wout[36][19] = 8'hAC;
    assign wout[36][20] = 8'hD0;
    assign wout[36][21] = 8'hF4;
    assign wout[36][22] = 8'h18;
    assign wout[36][23] = 8'h3C;
    assign wout[36][24] = 8'h60;
    assign wout[36][25] = 8'h84;
    assign wout[36][26] = 8'hA8;
    assign wout[36][27] = 8'hCC;
    assign wout[36][28] = 8'hF0;
    assign wout[36][29] = 8'h14;
    assign wout[36][30] = 8'h38;
    assign wout[36][31] = 8'h5C;
    assign wout[36][32] = 8'h80;
    assign wout[36][33] = 8'hA4;
    assign wout[36][34] = 8'hC8;
    assign wout[36][35] = 8'hEC;
    assign wout[36][36] = 8'h10;
    assign wout[36][37] = 8'h34;
    assign wout[36][38] = 8'h58;
    assign wout[36][39] = 8'h7C;
    assign wout[36][40] = 8'hA0;
    assign wout[36][41] = 8'hC4;
    assign wout[36][42] = 8'hE8;
    assign wout[36][43] = 8'h0C;
    assign wout[36][44] = 8'h30;
    assign wout[36][45] = 8'h54;
    assign wout[36][46] = 8'h78;
    assign wout[36][47] = 8'h9C;
    assign wout[36][48] = 8'hC0;
    assign wout[36][49] = 8'hE4;
    assign wout[36][50] = 8'h08;
    assign wout[36][51] = 8'h2C;
    assign wout[36][52] = 8'h50;
    assign wout[36][53] = 8'h74;
    assign wout[36][54] = 8'h98;
    assign wout[36][55] = 8'hBC;
    assign wout[36][56] = 8'hE0;
    assign wout[36][57] = 8'h04;
    assign wout[36][58] = 8'h28;
    assign wout[36][59] = 8'h4C;
    assign wout[36][60] = 8'h70;
    assign wout[36][61] = 8'h94;
    assign wout[36][62] = 8'hB8;
    assign wout[36][63] = 8'hDC;
    assign wout[37][0] = 8'h00;
    assign wout[37][1] = 8'h25;
    assign wout[37][2] = 8'h4A;
    assign wout[37][3] = 8'h6F;
    assign wout[37][4] = 8'h94;
    assign wout[37][5] = 8'hB9;
    assign wout[37][6] = 8'hDE;
    assign wout[37][7] = 8'h03;
    assign wout[37][8] = 8'h28;
    assign wout[37][9] = 8'h4D;
    assign wout[37][10] = 8'h72;
    assign wout[37][11] = 8'h97;
    assign wout[37][12] = 8'hBC;
    assign wout[37][13] = 8'hE1;
    assign wout[37][14] = 8'h06;
    assign wout[37][15] = 8'h2B;
    assign wout[37][16] = 8'h50;
    assign wout[37][17] = 8'h75;
    assign wout[37][18] = 8'h9A;
    assign wout[37][19] = 8'hBF;
    assign wout[37][20] = 8'hE4;
    assign wout[37][21] = 8'h09;
    assign wout[37][22] = 8'h2E;
    assign wout[37][23] = 8'h53;
    assign wout[37][24] = 8'h78;
    assign wout[37][25] = 8'h9D;
    assign wout[37][26] = 8'hC2;
    assign wout[37][27] = 8'hE7;
    assign wout[37][28] = 8'h0C;
    assign wout[37][29] = 8'h31;
    assign wout[37][30] = 8'h56;
    assign wout[37][31] = 8'h7B;
    assign wout[37][32] = 8'hA0;
    assign wout[37][33] = 8'hC5;
    assign wout[37][34] = 8'hEA;
    assign wout[37][35] = 8'h0F;
    assign wout[37][36] = 8'h34;
    assign wout[37][37] = 8'h59;
    assign wout[37][38] = 8'h7E;
    assign wout[37][39] = 8'hA3;
    assign wout[37][40] = 8'hC8;
    assign wout[37][41] = 8'hED;
    assign wout[37][42] = 8'h12;
    assign wout[37][43] = 8'h37;
    assign wout[37][44] = 8'h5C;
    assign wout[37][45] = 8'h81;
    assign wout[37][46] = 8'hA6;
    assign wout[37][47] = 8'hCB;
    assign wout[37][48] = 8'hF0;
    assign wout[37][49] = 8'h15;
    assign wout[37][50] = 8'h3A;
    assign wout[37][51] = 8'h5F;
    assign wout[37][52] = 8'h84;
    assign wout[37][53] = 8'hA9;
    assign wout[37][54] = 8'hCE;
    assign wout[37][55] = 8'hF3;
    assign wout[37][56] = 8'h18;
    assign wout[37][57] = 8'h3D;
    assign wout[37][58] = 8'h62;
    assign wout[37][59] = 8'h87;
    assign wout[37][60] = 8'hAC;
    assign wout[37][61] = 8'hD1;
    assign wout[37][62] = 8'hF6;
    assign wout[37][63] = 8'h1B;
    assign wout[38][0] = 8'h00;
    assign wout[38][1] = 8'h26;
    assign wout[38][2] = 8'h4C;
    assign wout[38][3] = 8'h72;
    assign wout[38][4] = 8'h98;
    assign wout[38][5] = 8'hBE;
    assign wout[38][6] = 8'hE4;
    assign wout[38][7] = 8'h0A;
    assign wout[38][8] = 8'h30;
    assign wout[38][9] = 8'h56;
    assign wout[38][10] = 8'h7C;
    assign wout[38][11] = 8'hA2;
    assign wout[38][12] = 8'hC8;
    assign wout[38][13] = 8'hEE;
    assign wout[38][14] = 8'h14;
    assign wout[38][15] = 8'h3A;
    assign wout[38][16] = 8'h60;
    assign wout[38][17] = 8'h86;
    assign wout[38][18] = 8'hAC;
    assign wout[38][19] = 8'hD2;
    assign wout[38][20] = 8'hF8;
    assign wout[38][21] = 8'h1E;
    assign wout[38][22] = 8'h44;
    assign wout[38][23] = 8'h6A;
    assign wout[38][24] = 8'h90;
    assign wout[38][25] = 8'hB6;
    assign wout[38][26] = 8'hDC;
    assign wout[38][27] = 8'h02;
    assign wout[38][28] = 8'h28;
    assign wout[38][29] = 8'h4E;
    assign wout[38][30] = 8'h74;
    assign wout[38][31] = 8'h9A;
    assign wout[38][32] = 8'hC0;
    assign wout[38][33] = 8'hE6;
    assign wout[38][34] = 8'h0C;
    assign wout[38][35] = 8'h32;
    assign wout[38][36] = 8'h58;
    assign wout[38][37] = 8'h7E;
    assign wout[38][38] = 8'hA4;
    assign wout[38][39] = 8'hCA;
    assign wout[38][40] = 8'hF0;
    assign wout[38][41] = 8'h16;
    assign wout[38][42] = 8'h3C;
    assign wout[38][43] = 8'h62;
    assign wout[38][44] = 8'h88;
    assign wout[38][45] = 8'hAE;
    assign wout[38][46] = 8'hD4;
    assign wout[38][47] = 8'hFA;
    assign wout[38][48] = 8'h20;
    assign wout[38][49] = 8'h46;
    assign wout[38][50] = 8'h6C;
    assign wout[38][51] = 8'h92;
    assign wout[38][52] = 8'hB8;
    assign wout[38][53] = 8'hDE;
    assign wout[38][54] = 8'h04;
    assign wout[38][55] = 8'h2A;
    assign wout[38][56] = 8'h50;
    assign wout[38][57] = 8'h76;
    assign wout[38][58] = 8'h9C;
    assign wout[38][59] = 8'hC2;
    assign wout[38][60] = 8'hE8;
    assign wout[38][61] = 8'h0E;
    assign wout[38][62] = 8'h34;
    assign wout[38][63] = 8'h5A;
    assign wout[39][0] = 8'h00;
    assign wout[39][1] = 8'h27;
    assign wout[39][2] = 8'h4E;
    assign wout[39][3] = 8'h75;
    assign wout[39][4] = 8'h9C;
    assign wout[39][5] = 8'hC3;
    assign wout[39][6] = 8'hEA;
    assign wout[39][7] = 8'h11;
    assign wout[39][8] = 8'h38;
    assign wout[39][9] = 8'h5F;
    assign wout[39][10] = 8'h86;
    assign wout[39][11] = 8'hAD;
    assign wout[39][12] = 8'hD4;
    assign wout[39][13] = 8'hFB;
    assign wout[39][14] = 8'h22;
    assign wout[39][15] = 8'h49;
    assign wout[39][16] = 8'h70;
    assign wout[39][17] = 8'h97;
    assign wout[39][18] = 8'hBE;
    assign wout[39][19] = 8'hE5;
    assign wout[39][20] = 8'h0C;
    assign wout[39][21] = 8'h33;
    assign wout[39][22] = 8'h5A;
    assign wout[39][23] = 8'h81;
    assign wout[39][24] = 8'hA8;
    assign wout[39][25] = 8'hCF;
    assign wout[39][26] = 8'hF6;
    assign wout[39][27] = 8'h1D;
    assign wout[39][28] = 8'h44;
    assign wout[39][29] = 8'h6B;
    assign wout[39][30] = 8'h92;
    assign wout[39][31] = 8'hB9;
    assign wout[39][32] = 8'hE0;
    assign wout[39][33] = 8'h07;
    assign wout[39][34] = 8'h2E;
    assign wout[39][35] = 8'h55;
    assign wout[39][36] = 8'h7C;
    assign wout[39][37] = 8'hA3;
    assign wout[39][38] = 8'hCA;
    assign wout[39][39] = 8'hF1;
    assign wout[39][40] = 8'h18;
    assign wout[39][41] = 8'h3F;
    assign wout[39][42] = 8'h66;
    assign wout[39][43] = 8'h8D;
    assign wout[39][44] = 8'hB4;
    assign wout[39][45] = 8'hDB;
    assign wout[39][46] = 8'h02;
    assign wout[39][47] = 8'h29;
    assign wout[39][48] = 8'h50;
    assign wout[39][49] = 8'h77;
    assign wout[39][50] = 8'h9E;
    assign wout[39][51] = 8'hC5;
    assign wout[39][52] = 8'hEC;
    assign wout[39][53] = 8'h13;
    assign wout[39][54] = 8'h3A;
    assign wout[39][55] = 8'h61;
    assign wout[39][56] = 8'h88;
    assign wout[39][57] = 8'hAF;
    assign wout[39][58] = 8'hD6;
    assign wout[39][59] = 8'hFD;
    assign wout[39][60] = 8'h24;
    assign wout[39][61] = 8'h4B;
    assign wout[39][62] = 8'h72;
    assign wout[39][63] = 8'h99;
    assign wout[40][0] = 8'h00;
    assign wout[40][1] = 8'h28;
    assign wout[40][2] = 8'h50;
    assign wout[40][3] = 8'h78;
    assign wout[40][4] = 8'hA0;
    assign wout[40][5] = 8'hC8;
    assign wout[40][6] = 8'hF0;
    assign wout[40][7] = 8'h18;
    assign wout[40][8] = 8'h40;
    assign wout[40][9] = 8'h68;
    assign wout[40][10] = 8'h90;
    assign wout[40][11] = 8'hB8;
    assign wout[40][12] = 8'hE0;
    assign wout[40][13] = 8'h08;
    assign wout[40][14] = 8'h30;
    assign wout[40][15] = 8'h58;
    assign wout[40][16] = 8'h80;
    assign wout[40][17] = 8'hA8;
    assign wout[40][18] = 8'hD0;
    assign wout[40][19] = 8'hF8;
    assign wout[40][20] = 8'h20;
    assign wout[40][21] = 8'h48;
    assign wout[40][22] = 8'h70;
    assign wout[40][23] = 8'h98;
    assign wout[40][24] = 8'hC0;
    assign wout[40][25] = 8'hE8;
    assign wout[40][26] = 8'h10;
    assign wout[40][27] = 8'h38;
    assign wout[40][28] = 8'h60;
    assign wout[40][29] = 8'h88;
    assign wout[40][30] = 8'hB0;
    assign wout[40][31] = 8'hD8;
    assign wout[40][32] = 8'h00;
    assign wout[40][33] = 8'h28;
    assign wout[40][34] = 8'h50;
    assign wout[40][35] = 8'h78;
    assign wout[40][36] = 8'hA0;
    assign wout[40][37] = 8'hC8;
    assign wout[40][38] = 8'hF0;
    assign wout[40][39] = 8'h18;
    assign wout[40][40] = 8'h40;
    assign wout[40][41] = 8'h68;
    assign wout[40][42] = 8'h90;
    assign wout[40][43] = 8'hB8;
    assign wout[40][44] = 8'hE0;
    assign wout[40][45] = 8'h08;
    assign wout[40][46] = 8'h30;
    assign wout[40][47] = 8'h58;
    assign wout[40][48] = 8'h80;
    assign wout[40][49] = 8'hA8;
    assign wout[40][50] = 8'hD0;
    assign wout[40][51] = 8'hF8;
    assign wout[40][52] = 8'h20;
    assign wout[40][53] = 8'h48;
    assign wout[40][54] = 8'h70;
    assign wout[40][55] = 8'h98;
    assign wout[40][56] = 8'hC0;
    assign wout[40][57] = 8'hE8;
    assign wout[40][58] = 8'h10;
    assign wout[40][59] = 8'h38;
    assign wout[40][60] = 8'h60;
    assign wout[40][61] = 8'h88;
    assign wout[40][62] = 8'hB0;
    assign wout[40][63] = 8'hD8;
    assign wout[41][0] = 8'h00;
    assign wout[41][1] = 8'h29;
    assign wout[41][2] = 8'h52;
    assign wout[41][3] = 8'h7B;
    assign wout[41][4] = 8'hA4;
    assign wout[41][5] = 8'hCD;
    assign wout[41][6] = 8'hF6;
    assign wout[41][7] = 8'h1F;
    assign wout[41][8] = 8'h48;
    assign wout[41][9] = 8'h71;
    assign wout[41][10] = 8'h9A;
    assign wout[41][11] = 8'hC3;
    assign wout[41][12] = 8'hEC;
    assign wout[41][13] = 8'h15;
    assign wout[41][14] = 8'h3E;
    assign wout[41][15] = 8'h67;
    assign wout[41][16] = 8'h90;
    assign wout[41][17] = 8'hB9;
    assign wout[41][18] = 8'hE2;
    assign wout[41][19] = 8'h0B;
    assign wout[41][20] = 8'h34;
    assign wout[41][21] = 8'h5D;
    assign wout[41][22] = 8'h86;
    assign wout[41][23] = 8'hAF;
    assign wout[41][24] = 8'hD8;
    assign wout[41][25] = 8'h01;
    assign wout[41][26] = 8'h2A;
    assign wout[41][27] = 8'h53;
    assign wout[41][28] = 8'h7C;
    assign wout[41][29] = 8'hA5;
    assign wout[41][30] = 8'hCE;
    assign wout[41][31] = 8'hF7;
    assign wout[41][32] = 8'h20;
    assign wout[41][33] = 8'h49;
    assign wout[41][34] = 8'h72;
    assign wout[41][35] = 8'h9B;
    assign wout[41][36] = 8'hC4;
    assign wout[41][37] = 8'hED;
    assign wout[41][38] = 8'h16;
    assign wout[41][39] = 8'h3F;
    assign wout[41][40] = 8'h68;
    assign wout[41][41] = 8'h91;
    assign wout[41][42] = 8'hBA;
    assign wout[41][43] = 8'hE3;
    assign wout[41][44] = 8'h0C;
    assign wout[41][45] = 8'h35;
    assign wout[41][46] = 8'h5E;
    assign wout[41][47] = 8'h87;
    assign wout[41][48] = 8'hB0;
    assign wout[41][49] = 8'hD9;
    assign wout[41][50] = 8'h02;
    assign wout[41][51] = 8'h2B;
    assign wout[41][52] = 8'h54;
    assign wout[41][53] = 8'h7D;
    assign wout[41][54] = 8'hA6;
    assign wout[41][55] = 8'hCF;
    assign wout[41][56] = 8'hF8;
    assign wout[41][57] = 8'h21;
    assign wout[41][58] = 8'h4A;
    assign wout[41][59] = 8'h73;
    assign wout[41][60] = 8'h9C;
    assign wout[41][61] = 8'hC5;
    assign wout[41][62] = 8'hEE;
    assign wout[41][63] = 8'h17;
    assign wout[42][0] = 8'h00;
    assign wout[42][1] = 8'h2A;
    assign wout[42][2] = 8'h54;
    assign wout[42][3] = 8'h7E;
    assign wout[42][4] = 8'hA8;
    assign wout[42][5] = 8'hD2;
    assign wout[42][6] = 8'hFC;
    assign wout[42][7] = 8'h26;
    assign wout[42][8] = 8'h50;
    assign wout[42][9] = 8'h7A;
    assign wout[42][10] = 8'hA4;
    assign wout[42][11] = 8'hCE;
    assign wout[42][12] = 8'hF8;
    assign wout[42][13] = 8'h22;
    assign wout[42][14] = 8'h4C;
    assign wout[42][15] = 8'h76;
    assign wout[42][16] = 8'hA0;
    assign wout[42][17] = 8'hCA;
    assign wout[42][18] = 8'hF4;
    assign wout[42][19] = 8'h1E;
    assign wout[42][20] = 8'h48;
    assign wout[42][21] = 8'h72;
    assign wout[42][22] = 8'h9C;
    assign wout[42][23] = 8'hC6;
    assign wout[42][24] = 8'hF0;
    assign wout[42][25] = 8'h1A;
    assign wout[42][26] = 8'h44;
    assign wout[42][27] = 8'h6E;
    assign wout[42][28] = 8'h98;
    assign wout[42][29] = 8'hC2;
    assign wout[42][30] = 8'hEC;
    assign wout[42][31] = 8'h16;
    assign wout[42][32] = 8'h40;
    assign wout[42][33] = 8'h6A;
    assign wout[42][34] = 8'h94;
    assign wout[42][35] = 8'hBE;
    assign wout[42][36] = 8'hE8;
    assign wout[42][37] = 8'h12;
    assign wout[42][38] = 8'h3C;
    assign wout[42][39] = 8'h66;
    assign wout[42][40] = 8'h90;
    assign wout[42][41] = 8'hBA;
    assign wout[42][42] = 8'hE4;
    assign wout[42][43] = 8'h0E;
    assign wout[42][44] = 8'h38;
    assign wout[42][45] = 8'h62;
    assign wout[42][46] = 8'h8C;
    assign wout[42][47] = 8'hB6;
    assign wout[42][48] = 8'hE0;
    assign wout[42][49] = 8'h0A;
    assign wout[42][50] = 8'h34;
    assign wout[42][51] = 8'h5E;
    assign wout[42][52] = 8'h88;
    assign wout[42][53] = 8'hB2;
    assign wout[42][54] = 8'hDC;
    assign wout[42][55] = 8'h06;
    assign wout[42][56] = 8'h30;
    assign wout[42][57] = 8'h5A;
    assign wout[42][58] = 8'h84;
    assign wout[42][59] = 8'hAE;
    assign wout[42][60] = 8'hD8;
    assign wout[42][61] = 8'h02;
    assign wout[42][62] = 8'h2C;
    assign wout[42][63] = 8'h56;
    assign wout[43][0] = 8'h00;
    assign wout[43][1] = 8'h2B;
    assign wout[43][2] = 8'h56;
    assign wout[43][3] = 8'h81;
    assign wout[43][4] = 8'hAC;
    assign wout[43][5] = 8'hD7;
    assign wout[43][6] = 8'h02;
    assign wout[43][7] = 8'h2D;
    assign wout[43][8] = 8'h58;
    assign wout[43][9] = 8'h83;
    assign wout[43][10] = 8'hAE;
    assign wout[43][11] = 8'hD9;
    assign wout[43][12] = 8'h04;
    assign wout[43][13] = 8'h2F;
    assign wout[43][14] = 8'h5A;
    assign wout[43][15] = 8'h85;
    assign wout[43][16] = 8'hB0;
    assign wout[43][17] = 8'hDB;
    assign wout[43][18] = 8'h06;
    assign wout[43][19] = 8'h31;
    assign wout[43][20] = 8'h5C;
    assign wout[43][21] = 8'h87;
    assign wout[43][22] = 8'hB2;
    assign wout[43][23] = 8'hDD;
    assign wout[43][24] = 8'h08;
    assign wout[43][25] = 8'h33;
    assign wout[43][26] = 8'h5E;
    assign wout[43][27] = 8'h89;
    assign wout[43][28] = 8'hB4;
    assign wout[43][29] = 8'hDF;
    assign wout[43][30] = 8'h0A;
    assign wout[43][31] = 8'h35;
    assign wout[43][32] = 8'h60;
    assign wout[43][33] = 8'h8B;
    assign wout[43][34] = 8'hB6;
    assign wout[43][35] = 8'hE1;
    assign wout[43][36] = 8'h0C;
    assign wout[43][37] = 8'h37;
    assign wout[43][38] = 8'h62;
    assign wout[43][39] = 8'h8D;
    assign wout[43][40] = 8'hB8;
    assign wout[43][41] = 8'hE3;
    assign wout[43][42] = 8'h0E;
    assign wout[43][43] = 8'h39;
    assign wout[43][44] = 8'h64;
    assign wout[43][45] = 8'h8F;
    assign wout[43][46] = 8'hBA;
    assign wout[43][47] = 8'hE5;
    assign wout[43][48] = 8'h10;
    assign wout[43][49] = 8'h3B;
    assign wout[43][50] = 8'h66;
    assign wout[43][51] = 8'h91;
    assign wout[43][52] = 8'hBC;
    assign wout[43][53] = 8'hE7;
    assign wout[43][54] = 8'h12;
    assign wout[43][55] = 8'h3D;
    assign wout[43][56] = 8'h68;
    assign wout[43][57] = 8'h93;
    assign wout[43][58] = 8'hBE;
    assign wout[43][59] = 8'hE9;
    assign wout[43][60] = 8'h14;
    assign wout[43][61] = 8'h3F;
    assign wout[43][62] = 8'h6A;
    assign wout[43][63] = 8'h95;
    assign wout[44][0] = 8'h00;
    assign wout[44][1] = 8'h2C;
    assign wout[44][2] = 8'h58;
    assign wout[44][3] = 8'h84;
    assign wout[44][4] = 8'hB0;
    assign wout[44][5] = 8'hDC;
    assign wout[44][6] = 8'h08;
    assign wout[44][7] = 8'h34;
    assign wout[44][8] = 8'h60;
    assign wout[44][9] = 8'h8C;
    assign wout[44][10] = 8'hB8;
    assign wout[44][11] = 8'hE4;
    assign wout[44][12] = 8'h10;
    assign wout[44][13] = 8'h3C;
    assign wout[44][14] = 8'h68;
    assign wout[44][15] = 8'h94;
    assign wout[44][16] = 8'hC0;
    assign wout[44][17] = 8'hEC;
    assign wout[44][18] = 8'h18;
    assign wout[44][19] = 8'h44;
    assign wout[44][20] = 8'h70;
    assign wout[44][21] = 8'h9C;
    assign wout[44][22] = 8'hC8;
    assign wout[44][23] = 8'hF4;
    assign wout[44][24] = 8'h20;
    assign wout[44][25] = 8'h4C;
    assign wout[44][26] = 8'h78;
    assign wout[44][27] = 8'hA4;
    assign wout[44][28] = 8'hD0;
    assign wout[44][29] = 8'hFC;
    assign wout[44][30] = 8'h28;
    assign wout[44][31] = 8'h54;
    assign wout[44][32] = 8'h80;
    assign wout[44][33] = 8'hAC;
    assign wout[44][34] = 8'hD8;
    assign wout[44][35] = 8'h04;
    assign wout[44][36] = 8'h30;
    assign wout[44][37] = 8'h5C;
    assign wout[44][38] = 8'h88;
    assign wout[44][39] = 8'hB4;
    assign wout[44][40] = 8'hE0;
    assign wout[44][41] = 8'h0C;
    assign wout[44][42] = 8'h38;
    assign wout[44][43] = 8'h64;
    assign wout[44][44] = 8'h90;
    assign wout[44][45] = 8'hBC;
    assign wout[44][46] = 8'hE8;
    assign wout[44][47] = 8'h14;
    assign wout[44][48] = 8'h40;
    assign wout[44][49] = 8'h6C;
    assign wout[44][50] = 8'h98;
    assign wout[44][51] = 8'hC4;
    assign wout[44][52] = 8'hF0;
    assign wout[44][53] = 8'h1C;
    assign wout[44][54] = 8'h48;
    assign wout[44][55] = 8'h74;
    assign wout[44][56] = 8'hA0;
    assign wout[44][57] = 8'hCC;
    assign wout[44][58] = 8'hF8;
    assign wout[44][59] = 8'h24;
    assign wout[44][60] = 8'h50;
    assign wout[44][61] = 8'h7C;
    assign wout[44][62] = 8'hA8;
    assign wout[44][63] = 8'hD4;
    assign wout[45][0] = 8'h00;
    assign wout[45][1] = 8'h2D;
    assign wout[45][2] = 8'h5A;
    assign wout[45][3] = 8'h87;
    assign wout[45][4] = 8'hB4;
    assign wout[45][5] = 8'hE1;
    assign wout[45][6] = 8'h0E;
    assign wout[45][7] = 8'h3B;
    assign wout[45][8] = 8'h68;
    assign wout[45][9] = 8'h95;
    assign wout[45][10] = 8'hC2;
    assign wout[45][11] = 8'hEF;
    assign wout[45][12] = 8'h1C;
    assign wout[45][13] = 8'h49;
    assign wout[45][14] = 8'h76;
    assign wout[45][15] = 8'hA3;
    assign wout[45][16] = 8'hD0;
    assign wout[45][17] = 8'hFD;
    assign wout[45][18] = 8'h2A;
    assign wout[45][19] = 8'h57;
    assign wout[45][20] = 8'h84;
    assign wout[45][21] = 8'hB1;
    assign wout[45][22] = 8'hDE;
    assign wout[45][23] = 8'h0B;
    assign wout[45][24] = 8'h38;
    assign wout[45][25] = 8'h65;
    assign wout[45][26] = 8'h92;
    assign wout[45][27] = 8'hBF;
    assign wout[45][28] = 8'hEC;
    assign wout[45][29] = 8'h19;
    assign wout[45][30] = 8'h46;
    assign wout[45][31] = 8'h73;
    assign wout[45][32] = 8'hA0;
    assign wout[45][33] = 8'hCD;
    assign wout[45][34] = 8'hFA;
    assign wout[45][35] = 8'h27;
    assign wout[45][36] = 8'h54;
    assign wout[45][37] = 8'h81;
    assign wout[45][38] = 8'hAE;
    assign wout[45][39] = 8'hDB;
    assign wout[45][40] = 8'h08;
    assign wout[45][41] = 8'h35;
    assign wout[45][42] = 8'h62;
    assign wout[45][43] = 8'h8F;
    assign wout[45][44] = 8'hBC;
    assign wout[45][45] = 8'hE9;
    assign wout[45][46] = 8'h16;
    assign wout[45][47] = 8'h43;
    assign wout[45][48] = 8'h70;
    assign wout[45][49] = 8'h9D;
    assign wout[45][50] = 8'hCA;
    assign wout[45][51] = 8'hF7;
    assign wout[45][52] = 8'h24;
    assign wout[45][53] = 8'h51;
    assign wout[45][54] = 8'h7E;
    assign wout[45][55] = 8'hAB;
    assign wout[45][56] = 8'hD8;
    assign wout[45][57] = 8'h05;
    assign wout[45][58] = 8'h32;
    assign wout[45][59] = 8'h5F;
    assign wout[45][60] = 8'h8C;
    assign wout[45][61] = 8'hB9;
    assign wout[45][62] = 8'hE6;
    assign wout[45][63] = 8'h13;
    assign wout[46][0] = 8'h00;
    assign wout[46][1] = 8'h2E;
    assign wout[46][2] = 8'h5C;
    assign wout[46][3] = 8'h8A;
    assign wout[46][4] = 8'hB8;
    assign wout[46][5] = 8'hE6;
    assign wout[46][6] = 8'h14;
    assign wout[46][7] = 8'h42;
    assign wout[46][8] = 8'h70;
    assign wout[46][9] = 8'h9E;
    assign wout[46][10] = 8'hCC;
    assign wout[46][11] = 8'hFA;
    assign wout[46][12] = 8'h28;
    assign wout[46][13] = 8'h56;
    assign wout[46][14] = 8'h84;
    assign wout[46][15] = 8'hB2;
    assign wout[46][16] = 8'hE0;
    assign wout[46][17] = 8'h0E;
    assign wout[46][18] = 8'h3C;
    assign wout[46][19] = 8'h6A;
    assign wout[46][20] = 8'h98;
    assign wout[46][21] = 8'hC6;
    assign wout[46][22] = 8'hF4;
    assign wout[46][23] = 8'h22;
    assign wout[46][24] = 8'h50;
    assign wout[46][25] = 8'h7E;
    assign wout[46][26] = 8'hAC;
    assign wout[46][27] = 8'hDA;
    assign wout[46][28] = 8'h08;
    assign wout[46][29] = 8'h36;
    assign wout[46][30] = 8'h64;
    assign wout[46][31] = 8'h92;
    assign wout[46][32] = 8'hC0;
    assign wout[46][33] = 8'hEE;
    assign wout[46][34] = 8'h1C;
    assign wout[46][35] = 8'h4A;
    assign wout[46][36] = 8'h78;
    assign wout[46][37] = 8'hA6;
    assign wout[46][38] = 8'hD4;
    assign wout[46][39] = 8'h02;
    assign wout[46][40] = 8'h30;
    assign wout[46][41] = 8'h5E;
    assign wout[46][42] = 8'h8C;
    assign wout[46][43] = 8'hBA;
    assign wout[46][44] = 8'hE8;
    assign wout[46][45] = 8'h16;
    assign wout[46][46] = 8'h44;
    assign wout[46][47] = 8'h72;
    assign wout[46][48] = 8'hA0;
    assign wout[46][49] = 8'hCE;
    assign wout[46][50] = 8'hFC;
    assign wout[46][51] = 8'h2A;
    assign wout[46][52] = 8'h58;
    assign wout[46][53] = 8'h86;
    assign wout[46][54] = 8'hB4;
    assign wout[46][55] = 8'hE2;
    assign wout[46][56] = 8'h10;
    assign wout[46][57] = 8'h3E;
    assign wout[46][58] = 8'h6C;
    assign wout[46][59] = 8'h9A;
    assign wout[46][60] = 8'hC8;
    assign wout[46][61] = 8'hF6;
    assign wout[46][62] = 8'h24;
    assign wout[46][63] = 8'h52;
    assign wout[47][0] = 8'h00;
    assign wout[47][1] = 8'h2F;
    assign wout[47][2] = 8'h5E;
    assign wout[47][3] = 8'h8D;
    assign wout[47][4] = 8'hBC;
    assign wout[47][5] = 8'hEB;
    assign wout[47][6] = 8'h1A;
    assign wout[47][7] = 8'h49;
    assign wout[47][8] = 8'h78;
    assign wout[47][9] = 8'hA7;
    assign wout[47][10] = 8'hD6;
    assign wout[47][11] = 8'h05;
    assign wout[47][12] = 8'h34;
    assign wout[47][13] = 8'h63;
    assign wout[47][14] = 8'h92;
    assign wout[47][15] = 8'hC1;
    assign wout[47][16] = 8'hF0;
    assign wout[47][17] = 8'h1F;
    assign wout[47][18] = 8'h4E;
    assign wout[47][19] = 8'h7D;
    assign wout[47][20] = 8'hAC;
    assign wout[47][21] = 8'hDB;
    assign wout[47][22] = 8'h0A;
    assign wout[47][23] = 8'h39;
    assign wout[47][24] = 8'h68;
    assign wout[47][25] = 8'h97;
    assign wout[47][26] = 8'hC6;
    assign wout[47][27] = 8'hF5;
    assign wout[47][28] = 8'h24;
    assign wout[47][29] = 8'h53;
    assign wout[47][30] = 8'h82;
    assign wout[47][31] = 8'hB1;
    assign wout[47][32] = 8'hE0;
    assign wout[47][33] = 8'h0F;
    assign wout[47][34] = 8'h3E;
    assign wout[47][35] = 8'h6D;
    assign wout[47][36] = 8'h9C;
    assign wout[47][37] = 8'hCB;
    assign wout[47][38] = 8'hFA;
    assign wout[47][39] = 8'h29;
    assign wout[47][40] = 8'h58;
    assign wout[47][41] = 8'h87;
    assign wout[47][42] = 8'hB6;
    assign wout[47][43] = 8'hE5;
    assign wout[47][44] = 8'h14;
    assign wout[47][45] = 8'h43;
    assign wout[47][46] = 8'h72;
    assign wout[47][47] = 8'hA1;
    assign wout[47][48] = 8'hD0;
    assign wout[47][49] = 8'hFF;
    assign wout[47][50] = 8'h2E;
    assign wout[47][51] = 8'h5D;
    assign wout[47][52] = 8'h8C;
    assign wout[47][53] = 8'hBB;
    assign wout[47][54] = 8'hEA;
    assign wout[47][55] = 8'h19;
    assign wout[47][56] = 8'h48;
    assign wout[47][57] = 8'h77;
    assign wout[47][58] = 8'hA6;
    assign wout[47][59] = 8'hD5;
    assign wout[47][60] = 8'h04;
    assign wout[47][61] = 8'h33;
    assign wout[47][62] = 8'h62;
    assign wout[47][63] = 8'h91;
    assign wout[48][0] = 8'h00;
    assign wout[48][1] = 8'h30;
    assign wout[48][2] = 8'h60;
    assign wout[48][3] = 8'h90;
    assign wout[48][4] = 8'hC0;
    assign wout[48][5] = 8'hF0;
    assign wout[48][6] = 8'h20;
    assign wout[48][7] = 8'h50;
    assign wout[48][8] = 8'h80;
    assign wout[48][9] = 8'hB0;
    assign wout[48][10] = 8'hE0;
    assign wout[48][11] = 8'h10;
    assign wout[48][12] = 8'h40;
    assign wout[48][13] = 8'h70;
    assign wout[48][14] = 8'hA0;
    assign wout[48][15] = 8'hD0;
    assign wout[48][16] = 8'h00;
    assign wout[48][17] = 8'h30;
    assign wout[48][18] = 8'h60;
    assign wout[48][19] = 8'h90;
    assign wout[48][20] = 8'hC0;
    assign wout[48][21] = 8'hF0;
    assign wout[48][22] = 8'h20;
    assign wout[48][23] = 8'h50;
    assign wout[48][24] = 8'h80;
    assign wout[48][25] = 8'hB0;
    assign wout[48][26] = 8'hE0;
    assign wout[48][27] = 8'h10;
    assign wout[48][28] = 8'h40;
    assign wout[48][29] = 8'h70;
    assign wout[48][30] = 8'hA0;
    assign wout[48][31] = 8'hD0;
    assign wout[48][32] = 8'h00;
    assign wout[48][33] = 8'h30;
    assign wout[48][34] = 8'h60;
    assign wout[48][35] = 8'h90;
    assign wout[48][36] = 8'hC0;
    assign wout[48][37] = 8'hF0;
    assign wout[48][38] = 8'h20;
    assign wout[48][39] = 8'h50;
    assign wout[48][40] = 8'h80;
    assign wout[48][41] = 8'hB0;
    assign wout[48][42] = 8'hE0;
    assign wout[48][43] = 8'h10;
    assign wout[48][44] = 8'h40;
    assign wout[48][45] = 8'h70;
    assign wout[48][46] = 8'hA0;
    assign wout[48][47] = 8'hD0;
    assign wout[48][48] = 8'h00;
    assign wout[48][49] = 8'h30;
    assign wout[48][50] = 8'h60;
    assign wout[48][51] = 8'h90;
    assign wout[48][52] = 8'hC0;
    assign wout[48][53] = 8'hF0;
    assign wout[48][54] = 8'h20;
    assign wout[48][55] = 8'h50;
    assign wout[48][56] = 8'h80;
    assign wout[48][57] = 8'hB0;
    assign wout[48][58] = 8'hE0;
    assign wout[48][59] = 8'h10;
    assign wout[48][60] = 8'h40;
    assign wout[48][61] = 8'h70;
    assign wout[48][62] = 8'hA0;
    assign wout[48][63] = 8'hD0;
    assign wout[49][0] = 8'h00;
    assign wout[49][1] = 8'h31;
    assign wout[49][2] = 8'h62;
    assign wout[49][3] = 8'h93;
    assign wout[49][4] = 8'hC4;
    assign wout[49][5] = 8'hF5;
    assign wout[49][6] = 8'h26;
    assign wout[49][7] = 8'h57;
    assign wout[49][8] = 8'h88;
    assign wout[49][9] = 8'hB9;
    assign wout[49][10] = 8'hEA;
    assign wout[49][11] = 8'h1B;
    assign wout[49][12] = 8'h4C;
    assign wout[49][13] = 8'h7D;
    assign wout[49][14] = 8'hAE;
    assign wout[49][15] = 8'hDF;
    assign wout[49][16] = 8'h10;
    assign wout[49][17] = 8'h41;
    assign wout[49][18] = 8'h72;
    assign wout[49][19] = 8'hA3;
    assign wout[49][20] = 8'hD4;
    assign wout[49][21] = 8'h05;
    assign wout[49][22] = 8'h36;
    assign wout[49][23] = 8'h67;
    assign wout[49][24] = 8'h98;
    assign wout[49][25] = 8'hC9;
    assign wout[49][26] = 8'hFA;
    assign wout[49][27] = 8'h2B;
    assign wout[49][28] = 8'h5C;
    assign wout[49][29] = 8'h8D;
    assign wout[49][30] = 8'hBE;
    assign wout[49][31] = 8'hEF;
    assign wout[49][32] = 8'h20;
    assign wout[49][33] = 8'h51;
    assign wout[49][34] = 8'h82;
    assign wout[49][35] = 8'hB3;
    assign wout[49][36] = 8'hE4;
    assign wout[49][37] = 8'h15;
    assign wout[49][38] = 8'h46;
    assign wout[49][39] = 8'h77;
    assign wout[49][40] = 8'hA8;
    assign wout[49][41] = 8'hD9;
    assign wout[49][42] = 8'h0A;
    assign wout[49][43] = 8'h3B;
    assign wout[49][44] = 8'h6C;
    assign wout[49][45] = 8'h9D;
    assign wout[49][46] = 8'hCE;
    assign wout[49][47] = 8'hFF;
    assign wout[49][48] = 8'h30;
    assign wout[49][49] = 8'h61;
    assign wout[49][50] = 8'h92;
    assign wout[49][51] = 8'hC3;
    assign wout[49][52] = 8'hF4;
    assign wout[49][53] = 8'h25;
    assign wout[49][54] = 8'h56;
    assign wout[49][55] = 8'h87;
    assign wout[49][56] = 8'hB8;
    assign wout[49][57] = 8'hE9;
    assign wout[49][58] = 8'h1A;
    assign wout[49][59] = 8'h4B;
    assign wout[49][60] = 8'h7C;
    assign wout[49][61] = 8'hAD;
    assign wout[49][62] = 8'hDE;
    assign wout[49][63] = 8'h0F;
    assign wout[50][0] = 8'h00;
    assign wout[50][1] = 8'h32;
    assign wout[50][2] = 8'h64;
    assign wout[50][3] = 8'h96;
    assign wout[50][4] = 8'hC8;
    assign wout[50][5] = 8'hFA;
    assign wout[50][6] = 8'h2C;
    assign wout[50][7] = 8'h5E;
    assign wout[50][8] = 8'h90;
    assign wout[50][9] = 8'hC2;
    assign wout[50][10] = 8'hF4;
    assign wout[50][11] = 8'h26;
    assign wout[50][12] = 8'h58;
    assign wout[50][13] = 8'h8A;
    assign wout[50][14] = 8'hBC;
    assign wout[50][15] = 8'hEE;
    assign wout[50][16] = 8'h20;
    assign wout[50][17] = 8'h52;
    assign wout[50][18] = 8'h84;
    assign wout[50][19] = 8'hB6;
    assign wout[50][20] = 8'hE8;
    assign wout[50][21] = 8'h1A;
    assign wout[50][22] = 8'h4C;
    assign wout[50][23] = 8'h7E;
    assign wout[50][24] = 8'hB0;
    assign wout[50][25] = 8'hE2;
    assign wout[50][26] = 8'h14;
    assign wout[50][27] = 8'h46;
    assign wout[50][28] = 8'h78;
    assign wout[50][29] = 8'hAA;
    assign wout[50][30] = 8'hDC;
    assign wout[50][31] = 8'h0E;
    assign wout[50][32] = 8'h40;
    assign wout[50][33] = 8'h72;
    assign wout[50][34] = 8'hA4;
    assign wout[50][35] = 8'hD6;
    assign wout[50][36] = 8'h08;
    assign wout[50][37] = 8'h3A;
    assign wout[50][38] = 8'h6C;
    assign wout[50][39] = 8'h9E;
    assign wout[50][40] = 8'hD0;
    assign wout[50][41] = 8'h02;
    assign wout[50][42] = 8'h34;
    assign wout[50][43] = 8'h66;
    assign wout[50][44] = 8'h98;
    assign wout[50][45] = 8'hCA;
    assign wout[50][46] = 8'hFC;
    assign wout[50][47] = 8'h2E;
    assign wout[50][48] = 8'h60;
    assign wout[50][49] = 8'h92;
    assign wout[50][50] = 8'hC4;
    assign wout[50][51] = 8'hF6;
    assign wout[50][52] = 8'h28;
    assign wout[50][53] = 8'h5A;
    assign wout[50][54] = 8'h8C;
    assign wout[50][55] = 8'hBE;
    assign wout[50][56] = 8'hF0;
    assign wout[50][57] = 8'h22;
    assign wout[50][58] = 8'h54;
    assign wout[50][59] = 8'h86;
    assign wout[50][60] = 8'hB8;
    assign wout[50][61] = 8'hEA;
    assign wout[50][62] = 8'h1C;
    assign wout[50][63] = 8'h4E;
    assign wout[51][0] = 8'h00;
    assign wout[51][1] = 8'h33;
    assign wout[51][2] = 8'h66;
    assign wout[51][3] = 8'h99;
    assign wout[51][4] = 8'hCC;
    assign wout[51][5] = 8'hFF;
    assign wout[51][6] = 8'h32;
    assign wout[51][7] = 8'h65;
    assign wout[51][8] = 8'h98;
    assign wout[51][9] = 8'hCB;
    assign wout[51][10] = 8'hFE;
    assign wout[51][11] = 8'h31;
    assign wout[51][12] = 8'h64;
    assign wout[51][13] = 8'h97;
    assign wout[51][14] = 8'hCA;
    assign wout[51][15] = 8'hFD;
    assign wout[51][16] = 8'h30;
    assign wout[51][17] = 8'h63;
    assign wout[51][18] = 8'h96;
    assign wout[51][19] = 8'hC9;
    assign wout[51][20] = 8'hFC;
    assign wout[51][21] = 8'h2F;
    assign wout[51][22] = 8'h62;
    assign wout[51][23] = 8'h95;
    assign wout[51][24] = 8'hC8;
    assign wout[51][25] = 8'hFB;
    assign wout[51][26] = 8'h2E;
    assign wout[51][27] = 8'h61;
    assign wout[51][28] = 8'h94;
    assign wout[51][29] = 8'hC7;
    assign wout[51][30] = 8'hFA;
    assign wout[51][31] = 8'h2D;
    assign wout[51][32] = 8'h60;
    assign wout[51][33] = 8'h93;
    assign wout[51][34] = 8'hC6;
    assign wout[51][35] = 8'hF9;
    assign wout[51][36] = 8'h2C;
    assign wout[51][37] = 8'h5F;
    assign wout[51][38] = 8'h92;
    assign wout[51][39] = 8'hC5;
    assign wout[51][40] = 8'hF8;
    assign wout[51][41] = 8'h2B;
    assign wout[51][42] = 8'h5E;
    assign wout[51][43] = 8'h91;
    assign wout[51][44] = 8'hC4;
    assign wout[51][45] = 8'hF7;
    assign wout[51][46] = 8'h2A;
    assign wout[51][47] = 8'h5D;
    assign wout[51][48] = 8'h90;
    assign wout[51][49] = 8'hC3;
    assign wout[51][50] = 8'hF6;
    assign wout[51][51] = 8'h29;
    assign wout[51][52] = 8'h5C;
    assign wout[51][53] = 8'h8F;
    assign wout[51][54] = 8'hC2;
    assign wout[51][55] = 8'hF5;
    assign wout[51][56] = 8'h28;
    assign wout[51][57] = 8'h5B;
    assign wout[51][58] = 8'h8E;
    assign wout[51][59] = 8'hC1;
    assign wout[51][60] = 8'hF4;
    assign wout[51][61] = 8'h27;
    assign wout[51][62] = 8'h5A;
    assign wout[51][63] = 8'h8D;
    assign wout[52][0] = 8'h00;
    assign wout[52][1] = 8'h34;
    assign wout[52][2] = 8'h68;
    assign wout[52][3] = 8'h9C;
    assign wout[52][4] = 8'hD0;
    assign wout[52][5] = 8'h04;
    assign wout[52][6] = 8'h38;
    assign wout[52][7] = 8'h6C;
    assign wout[52][8] = 8'hA0;
    assign wout[52][9] = 8'hD4;
    assign wout[52][10] = 8'h08;
    assign wout[52][11] = 8'h3C;
    assign wout[52][12] = 8'h70;
    assign wout[52][13] = 8'hA4;
    assign wout[52][14] = 8'hD8;
    assign wout[52][15] = 8'h0C;
    assign wout[52][16] = 8'h40;
    assign wout[52][17] = 8'h74;
    assign wout[52][18] = 8'hA8;
    assign wout[52][19] = 8'hDC;
    assign wout[52][20] = 8'h10;
    assign wout[52][21] = 8'h44;
    assign wout[52][22] = 8'h78;
    assign wout[52][23] = 8'hAC;
    assign wout[52][24] = 8'hE0;
    assign wout[52][25] = 8'h14;
    assign wout[52][26] = 8'h48;
    assign wout[52][27] = 8'h7C;
    assign wout[52][28] = 8'hB0;
    assign wout[52][29] = 8'hE4;
    assign wout[52][30] = 8'h18;
    assign wout[52][31] = 8'h4C;
    assign wout[52][32] = 8'h80;
    assign wout[52][33] = 8'hB4;
    assign wout[52][34] = 8'hE8;
    assign wout[52][35] = 8'h1C;
    assign wout[52][36] = 8'h50;
    assign wout[52][37] = 8'h84;
    assign wout[52][38] = 8'hB8;
    assign wout[52][39] = 8'hEC;
    assign wout[52][40] = 8'h20;
    assign wout[52][41] = 8'h54;
    assign wout[52][42] = 8'h88;
    assign wout[52][43] = 8'hBC;
    assign wout[52][44] = 8'hF0;
    assign wout[52][45] = 8'h24;
    assign wout[52][46] = 8'h58;
    assign wout[52][47] = 8'h8C;
    assign wout[52][48] = 8'hC0;
    assign wout[52][49] = 8'hF4;
    assign wout[52][50] = 8'h28;
    assign wout[52][51] = 8'h5C;
    assign wout[52][52] = 8'h90;
    assign wout[52][53] = 8'hC4;
    assign wout[52][54] = 8'hF8;
    assign wout[52][55] = 8'h2C;
    assign wout[52][56] = 8'h60;
    assign wout[52][57] = 8'h94;
    assign wout[52][58] = 8'hC8;
    assign wout[52][59] = 8'hFC;
    assign wout[52][60] = 8'h30;
    assign wout[52][61] = 8'h64;
    assign wout[52][62] = 8'h98;
    assign wout[52][63] = 8'hCC;
    assign wout[53][0] = 8'h00;
    assign wout[53][1] = 8'h35;
    assign wout[53][2] = 8'h6A;
    assign wout[53][3] = 8'h9F;
    assign wout[53][4] = 8'hD4;
    assign wout[53][5] = 8'h09;
    assign wout[53][6] = 8'h3E;
    assign wout[53][7] = 8'h73;
    assign wout[53][8] = 8'hA8;
    assign wout[53][9] = 8'hDD;
    assign wout[53][10] = 8'h12;
    assign wout[53][11] = 8'h47;
    assign wout[53][12] = 8'h7C;
    assign wout[53][13] = 8'hB1;
    assign wout[53][14] = 8'hE6;
    assign wout[53][15] = 8'h1B;
    assign wout[53][16] = 8'h50;
    assign wout[53][17] = 8'h85;
    assign wout[53][18] = 8'hBA;
    assign wout[53][19] = 8'hEF;
    assign wout[53][20] = 8'h24;
    assign wout[53][21] = 8'h59;
    assign wout[53][22] = 8'h8E;
    assign wout[53][23] = 8'hC3;
    assign wout[53][24] = 8'hF8;
    assign wout[53][25] = 8'h2D;
    assign wout[53][26] = 8'h62;
    assign wout[53][27] = 8'h97;
    assign wout[53][28] = 8'hCC;
    assign wout[53][29] = 8'h01;
    assign wout[53][30] = 8'h36;
    assign wout[53][31] = 8'h6B;
    assign wout[53][32] = 8'hA0;
    assign wout[53][33] = 8'hD5;
    assign wout[53][34] = 8'h0A;
    assign wout[53][35] = 8'h3F;
    assign wout[53][36] = 8'h74;
    assign wout[53][37] = 8'hA9;
    assign wout[53][38] = 8'hDE;
    assign wout[53][39] = 8'h13;
    assign wout[53][40] = 8'h48;
    assign wout[53][41] = 8'h7D;
    assign wout[53][42] = 8'hB2;
    assign wout[53][43] = 8'hE7;
    assign wout[53][44] = 8'h1C;
    assign wout[53][45] = 8'h51;
    assign wout[53][46] = 8'h86;
    assign wout[53][47] = 8'hBB;
    assign wout[53][48] = 8'hF0;
    assign wout[53][49] = 8'h25;
    assign wout[53][50] = 8'h5A;
    assign wout[53][51] = 8'h8F;
    assign wout[53][52] = 8'hC4;
    assign wout[53][53] = 8'hF9;
    assign wout[53][54] = 8'h2E;
    assign wout[53][55] = 8'h63;
    assign wout[53][56] = 8'h98;
    assign wout[53][57] = 8'hCD;
    assign wout[53][58] = 8'h02;
    assign wout[53][59] = 8'h37;
    assign wout[53][60] = 8'h6C;
    assign wout[53][61] = 8'hA1;
    assign wout[53][62] = 8'hD6;
    assign wout[53][63] = 8'h0B;
    assign wout[54][0] = 8'h00;
    assign wout[54][1] = 8'h36;
    assign wout[54][2] = 8'h6C;
    assign wout[54][3] = 8'hA2;
    assign wout[54][4] = 8'hD8;
    assign wout[54][5] = 8'h0E;
    assign wout[54][6] = 8'h44;
    assign wout[54][7] = 8'h7A;
    assign wout[54][8] = 8'hB0;
    assign wout[54][9] = 8'hE6;
    assign wout[54][10] = 8'h1C;
    assign wout[54][11] = 8'h52;
    assign wout[54][12] = 8'h88;
    assign wout[54][13] = 8'hBE;
    assign wout[54][14] = 8'hF4;
    assign wout[54][15] = 8'h2A;
    assign wout[54][16] = 8'h60;
    assign wout[54][17] = 8'h96;
    assign wout[54][18] = 8'hCC;
    assign wout[54][19] = 8'h02;
    assign wout[54][20] = 8'h38;
    assign wout[54][21] = 8'h6E;
    assign wout[54][22] = 8'hA4;
    assign wout[54][23] = 8'hDA;
    assign wout[54][24] = 8'h10;
    assign wout[54][25] = 8'h46;
    assign wout[54][26] = 8'h7C;
    assign wout[54][27] = 8'hB2;
    assign wout[54][28] = 8'hE8;
    assign wout[54][29] = 8'h1E;
    assign wout[54][30] = 8'h54;
    assign wout[54][31] = 8'h8A;
    assign wout[54][32] = 8'hC0;
    assign wout[54][33] = 8'hF6;
    assign wout[54][34] = 8'h2C;
    assign wout[54][35] = 8'h62;
    assign wout[54][36] = 8'h98;
    assign wout[54][37] = 8'hCE;
    assign wout[54][38] = 8'h04;
    assign wout[54][39] = 8'h3A;
    assign wout[54][40] = 8'h70;
    assign wout[54][41] = 8'hA6;
    assign wout[54][42] = 8'hDC;
    assign wout[54][43] = 8'h12;
    assign wout[54][44] = 8'h48;
    assign wout[54][45] = 8'h7E;
    assign wout[54][46] = 8'hB4;
    assign wout[54][47] = 8'hEA;
    assign wout[54][48] = 8'h20;
    assign wout[54][49] = 8'h56;
    assign wout[54][50] = 8'h8C;
    assign wout[54][51] = 8'hC2;
    assign wout[54][52] = 8'hF8;
    assign wout[54][53] = 8'h2E;
    assign wout[54][54] = 8'h64;
    assign wout[54][55] = 8'h9A;
    assign wout[54][56] = 8'hD0;
    assign wout[54][57] = 8'h06;
    assign wout[54][58] = 8'h3C;
    assign wout[54][59] = 8'h72;
    assign wout[54][60] = 8'hA8;
    assign wout[54][61] = 8'hDE;
    assign wout[54][62] = 8'h14;
    assign wout[54][63] = 8'h4A;
    assign wout[55][0] = 8'h00;
    assign wout[55][1] = 8'h37;
    assign wout[55][2] = 8'h6E;
    assign wout[55][3] = 8'hA5;
    assign wout[55][4] = 8'hDC;
    assign wout[55][5] = 8'h13;
    assign wout[55][6] = 8'h4A;
    assign wout[55][7] = 8'h81;
    assign wout[55][8] = 8'hB8;
    assign wout[55][9] = 8'hEF;
    assign wout[55][10] = 8'h26;
    assign wout[55][11] = 8'h5D;
    assign wout[55][12] = 8'h94;
    assign wout[55][13] = 8'hCB;
    assign wout[55][14] = 8'h02;
    assign wout[55][15] = 8'h39;
    assign wout[55][16] = 8'h70;
    assign wout[55][17] = 8'hA7;
    assign wout[55][18] = 8'hDE;
    assign wout[55][19] = 8'h15;
    assign wout[55][20] = 8'h4C;
    assign wout[55][21] = 8'h83;
    assign wout[55][22] = 8'hBA;
    assign wout[55][23] = 8'hF1;
    assign wout[55][24] = 8'h28;
    assign wout[55][25] = 8'h5F;
    assign wout[55][26] = 8'h96;
    assign wout[55][27] = 8'hCD;
    assign wout[55][28] = 8'h04;
    assign wout[55][29] = 8'h3B;
    assign wout[55][30] = 8'h72;
    assign wout[55][31] = 8'hA9;
    assign wout[55][32] = 8'hE0;
    assign wout[55][33] = 8'h17;
    assign wout[55][34] = 8'h4E;
    assign wout[55][35] = 8'h85;
    assign wout[55][36] = 8'hBC;
    assign wout[55][37] = 8'hF3;
    assign wout[55][38] = 8'h2A;
    assign wout[55][39] = 8'h61;
    assign wout[55][40] = 8'h98;
    assign wout[55][41] = 8'hCF;
    assign wout[55][42] = 8'h06;
    assign wout[55][43] = 8'h3D;
    assign wout[55][44] = 8'h74;
    assign wout[55][45] = 8'hAB;
    assign wout[55][46] = 8'hE2;
    assign wout[55][47] = 8'h19;
    assign wout[55][48] = 8'h50;
    assign wout[55][49] = 8'h87;
    assign wout[55][50] = 8'hBE;
    assign wout[55][51] = 8'hF5;
    assign wout[55][52] = 8'h2C;
    assign wout[55][53] = 8'h63;
    assign wout[55][54] = 8'h9A;
    assign wout[55][55] = 8'hD1;
    assign wout[55][56] = 8'h08;
    assign wout[55][57] = 8'h3F;
    assign wout[55][58] = 8'h76;
    assign wout[55][59] = 8'hAD;
    assign wout[55][60] = 8'hE4;
    assign wout[55][61] = 8'h1B;
    assign wout[55][62] = 8'h52;
    assign wout[55][63] = 8'h89;
    assign wout[56][0] = 8'h00;
    assign wout[56][1] = 8'h38;
    assign wout[56][2] = 8'h70;
    assign wout[56][3] = 8'hA8;
    assign wout[56][4] = 8'hE0;
    assign wout[56][5] = 8'h18;
    assign wout[56][6] = 8'h50;
    assign wout[56][7] = 8'h88;
    assign wout[56][8] = 8'hC0;
    assign wout[56][9] = 8'hF8;
    assign wout[56][10] = 8'h30;
    assign wout[56][11] = 8'h68;
    assign wout[56][12] = 8'hA0;
    assign wout[56][13] = 8'hD8;
    assign wout[56][14] = 8'h10;
    assign wout[56][15] = 8'h48;
    assign wout[56][16] = 8'h80;
    assign wout[56][17] = 8'hB8;
    assign wout[56][18] = 8'hF0;
    assign wout[56][19] = 8'h28;
    assign wout[56][20] = 8'h60;
    assign wout[56][21] = 8'h98;
    assign wout[56][22] = 8'hD0;
    assign wout[56][23] = 8'h08;
    assign wout[56][24] = 8'h40;
    assign wout[56][25] = 8'h78;
    assign wout[56][26] = 8'hB0;
    assign wout[56][27] = 8'hE8;
    assign wout[56][28] = 8'h20;
    assign wout[56][29] = 8'h58;
    assign wout[56][30] = 8'h90;
    assign wout[56][31] = 8'hC8;
    assign wout[56][32] = 8'h00;
    assign wout[56][33] = 8'h38;
    assign wout[56][34] = 8'h70;
    assign wout[56][35] = 8'hA8;
    assign wout[56][36] = 8'hE0;
    assign wout[56][37] = 8'h18;
    assign wout[56][38] = 8'h50;
    assign wout[56][39] = 8'h88;
    assign wout[56][40] = 8'hC0;
    assign wout[56][41] = 8'hF8;
    assign wout[56][42] = 8'h30;
    assign wout[56][43] = 8'h68;
    assign wout[56][44] = 8'hA0;
    assign wout[56][45] = 8'hD8;
    assign wout[56][46] = 8'h10;
    assign wout[56][47] = 8'h48;
    assign wout[56][48] = 8'h80;
    assign wout[56][49] = 8'hB8;
    assign wout[56][50] = 8'hF0;
    assign wout[56][51] = 8'h28;
    assign wout[56][52] = 8'h60;
    assign wout[56][53] = 8'h98;
    assign wout[56][54] = 8'hD0;
    assign wout[56][55] = 8'h08;
    assign wout[56][56] = 8'h40;
    assign wout[56][57] = 8'h78;
    assign wout[56][58] = 8'hB0;
    assign wout[56][59] = 8'hE8;
    assign wout[56][60] = 8'h20;
    assign wout[56][61] = 8'h58;
    assign wout[56][62] = 8'h90;
    assign wout[56][63] = 8'hC8;
    assign wout[57][0] = 8'h00;
    assign wout[57][1] = 8'h39;
    assign wout[57][2] = 8'h72;
    assign wout[57][3] = 8'hAB;
    assign wout[57][4] = 8'hE4;
    assign wout[57][5] = 8'h1D;
    assign wout[57][6] = 8'h56;
    assign wout[57][7] = 8'h8F;
    assign wout[57][8] = 8'hC8;
    assign wout[57][9] = 8'h01;
    assign wout[57][10] = 8'h3A;
    assign wout[57][11] = 8'h73;
    assign wout[57][12] = 8'hAC;
    assign wout[57][13] = 8'hE5;
    assign wout[57][14] = 8'h1E;
    assign wout[57][15] = 8'h57;
    assign wout[57][16] = 8'h90;
    assign wout[57][17] = 8'hC9;
    assign wout[57][18] = 8'h02;
    assign wout[57][19] = 8'h3B;
    assign wout[57][20] = 8'h74;
    assign wout[57][21] = 8'hAD;
    assign wout[57][22] = 8'hE6;
    assign wout[57][23] = 8'h1F;
    assign wout[57][24] = 8'h58;
    assign wout[57][25] = 8'h91;
    assign wout[57][26] = 8'hCA;
    assign wout[57][27] = 8'h03;
    assign wout[57][28] = 8'h3C;
    assign wout[57][29] = 8'h75;
    assign wout[57][30] = 8'hAE;
    assign wout[57][31] = 8'hE7;
    assign wout[57][32] = 8'h20;
    assign wout[57][33] = 8'h59;
    assign wout[57][34] = 8'h92;
    assign wout[57][35] = 8'hCB;
    assign wout[57][36] = 8'h04;
    assign wout[57][37] = 8'h3D;
    assign wout[57][38] = 8'h76;
    assign wout[57][39] = 8'hAF;
    assign wout[57][40] = 8'hE8;
    assign wout[57][41] = 8'h21;
    assign wout[57][42] = 8'h5A;
    assign wout[57][43] = 8'h93;
    assign wout[57][44] = 8'hCC;
    assign wout[57][45] = 8'h05;
    assign wout[57][46] = 8'h3E;
    assign wout[57][47] = 8'h77;
    assign wout[57][48] = 8'hB0;
    assign wout[57][49] = 8'hE9;
    assign wout[57][50] = 8'h22;
    assign wout[57][51] = 8'h5B;
    assign wout[57][52] = 8'h94;
    assign wout[57][53] = 8'hCD;
    assign wout[57][54] = 8'h06;
    assign wout[57][55] = 8'h3F;
    assign wout[57][56] = 8'h78;
    assign wout[57][57] = 8'hB1;
    assign wout[57][58] = 8'hEA;
    assign wout[57][59] = 8'h23;
    assign wout[57][60] = 8'h5C;
    assign wout[57][61] = 8'h95;
    assign wout[57][62] = 8'hCE;
    assign wout[57][63] = 8'h07;
    assign wout[58][0] = 8'h00;
    assign wout[58][1] = 8'h3A;
    assign wout[58][2] = 8'h74;
    assign wout[58][3] = 8'hAE;
    assign wout[58][4] = 8'hE8;
    assign wout[58][5] = 8'h22;
    assign wout[58][6] = 8'h5C;
    assign wout[58][7] = 8'h96;
    assign wout[58][8] = 8'hD0;
    assign wout[58][9] = 8'h0A;
    assign wout[58][10] = 8'h44;
    assign wout[58][11] = 8'h7E;
    assign wout[58][12] = 8'hB8;
    assign wout[58][13] = 8'hF2;
    assign wout[58][14] = 8'h2C;
    assign wout[58][15] = 8'h66;
    assign wout[58][16] = 8'hA0;
    assign wout[58][17] = 8'hDA;
    assign wout[58][18] = 8'h14;
    assign wout[58][19] = 8'h4E;
    assign wout[58][20] = 8'h88;
    assign wout[58][21] = 8'hC2;
    assign wout[58][22] = 8'hFC;
    assign wout[58][23] = 8'h36;
    assign wout[58][24] = 8'h70;
    assign wout[58][25] = 8'hAA;
    assign wout[58][26] = 8'hE4;
    assign wout[58][27] = 8'h1E;
    assign wout[58][28] = 8'h58;
    assign wout[58][29] = 8'h92;
    assign wout[58][30] = 8'hCC;
    assign wout[58][31] = 8'h06;
    assign wout[58][32] = 8'h40;
    assign wout[58][33] = 8'h7A;
    assign wout[58][34] = 8'hB4;
    assign wout[58][35] = 8'hEE;
    assign wout[58][36] = 8'h28;
    assign wout[58][37] = 8'h62;
    assign wout[58][38] = 8'h9C;
    assign wout[58][39] = 8'hD6;
    assign wout[58][40] = 8'h10;
    assign wout[58][41] = 8'h4A;
    assign wout[58][42] = 8'h84;
    assign wout[58][43] = 8'hBE;
    assign wout[58][44] = 8'hF8;
    assign wout[58][45] = 8'h32;
    assign wout[58][46] = 8'h6C;
    assign wout[58][47] = 8'hA6;
    assign wout[58][48] = 8'hE0;
    assign wout[58][49] = 8'h1A;
    assign wout[58][50] = 8'h54;
    assign wout[58][51] = 8'h8E;
    assign wout[58][52] = 8'hC8;
    assign wout[58][53] = 8'h02;
    assign wout[58][54] = 8'h3C;
    assign wout[58][55] = 8'h76;
    assign wout[58][56] = 8'hB0;
    assign wout[58][57] = 8'hEA;
    assign wout[58][58] = 8'h24;
    assign wout[58][59] = 8'h5E;
    assign wout[58][60] = 8'h98;
    assign wout[58][61] = 8'hD2;
    assign wout[58][62] = 8'h0C;
    assign wout[58][63] = 8'h46;
    assign wout[59][0] = 8'h00;
    assign wout[59][1] = 8'h3B;
    assign wout[59][2] = 8'h76;
    assign wout[59][3] = 8'hB1;
    assign wout[59][4] = 8'hEC;
    assign wout[59][5] = 8'h27;
    assign wout[59][6] = 8'h62;
    assign wout[59][7] = 8'h9D;
    assign wout[59][8] = 8'hD8;
    assign wout[59][9] = 8'h13;
    assign wout[59][10] = 8'h4E;
    assign wout[59][11] = 8'h89;
    assign wout[59][12] = 8'hC4;
    assign wout[59][13] = 8'hFF;
    assign wout[59][14] = 8'h3A;
    assign wout[59][15] = 8'h75;
    assign wout[59][16] = 8'hB0;
    assign wout[59][17] = 8'hEB;
    assign wout[59][18] = 8'h26;
    assign wout[59][19] = 8'h61;
    assign wout[59][20] = 8'h9C;
    assign wout[59][21] = 8'hD7;
    assign wout[59][22] = 8'h12;
    assign wout[59][23] = 8'h4D;
    assign wout[59][24] = 8'h88;
    assign wout[59][25] = 8'hC3;
    assign wout[59][26] = 8'hFE;
    assign wout[59][27] = 8'h39;
    assign wout[59][28] = 8'h74;
    assign wout[59][29] = 8'hAF;
    assign wout[59][30] = 8'hEA;
    assign wout[59][31] = 8'h25;
    assign wout[59][32] = 8'h60;
    assign wout[59][33] = 8'h9B;
    assign wout[59][34] = 8'hD6;
    assign wout[59][35] = 8'h11;
    assign wout[59][36] = 8'h4C;
    assign wout[59][37] = 8'h87;
    assign wout[59][38] = 8'hC2;
    assign wout[59][39] = 8'hFD;
    assign wout[59][40] = 8'h38;
    assign wout[59][41] = 8'h73;
    assign wout[59][42] = 8'hAE;
    assign wout[59][43] = 8'hE9;
    assign wout[59][44] = 8'h24;
    assign wout[59][45] = 8'h5F;
    assign wout[59][46] = 8'h9A;
    assign wout[59][47] = 8'hD5;
    assign wout[59][48] = 8'h10;
    assign wout[59][49] = 8'h4B;
    assign wout[59][50] = 8'h86;
    assign wout[59][51] = 8'hC1;
    assign wout[59][52] = 8'hFC;
    assign wout[59][53] = 8'h37;
    assign wout[59][54] = 8'h72;
    assign wout[59][55] = 8'hAD;
    assign wout[59][56] = 8'hE8;
    assign wout[59][57] = 8'h23;
    assign wout[59][58] = 8'h5E;
    assign wout[59][59] = 8'h99;
    assign wout[59][60] = 8'hD4;
    assign wout[59][61] = 8'h0F;
    assign wout[59][62] = 8'h4A;
    assign wout[59][63] = 8'h85;
    assign wout[60][0] = 8'h00;
    assign wout[60][1] = 8'h3C;
    assign wout[60][2] = 8'h78;
    assign wout[60][3] = 8'hB4;
    assign wout[60][4] = 8'hF0;
    assign wout[60][5] = 8'h2C;
    assign wout[60][6] = 8'h68;
    assign wout[60][7] = 8'hA4;
    assign wout[60][8] = 8'hE0;
    assign wout[60][9] = 8'h1C;
    assign wout[60][10] = 8'h58;
    assign wout[60][11] = 8'h94;
    assign wout[60][12] = 8'hD0;
    assign wout[60][13] = 8'h0C;
    assign wout[60][14] = 8'h48;
    assign wout[60][15] = 8'h84;
    assign wout[60][16] = 8'hC0;
    assign wout[60][17] = 8'hFC;
    assign wout[60][18] = 8'h38;
    assign wout[60][19] = 8'h74;
    assign wout[60][20] = 8'hB0;
    assign wout[60][21] = 8'hEC;
    assign wout[60][22] = 8'h28;
    assign wout[60][23] = 8'h64;
    assign wout[60][24] = 8'hA0;
    assign wout[60][25] = 8'hDC;
    assign wout[60][26] = 8'h18;
    assign wout[60][27] = 8'h54;
    assign wout[60][28] = 8'h90;
    assign wout[60][29] = 8'hCC;
    assign wout[60][30] = 8'h08;
    assign wout[60][31] = 8'h44;
    assign wout[60][32] = 8'h80;
    assign wout[60][33] = 8'hBC;
    assign wout[60][34] = 8'hF8;
    assign wout[60][35] = 8'h34;
    assign wout[60][36] = 8'h70;
    assign wout[60][37] = 8'hAC;
    assign wout[60][38] = 8'hE8;
    assign wout[60][39] = 8'h24;
    assign wout[60][40] = 8'h60;
    assign wout[60][41] = 8'h9C;
    assign wout[60][42] = 8'hD8;
    assign wout[60][43] = 8'h14;
    assign wout[60][44] = 8'h50;
    assign wout[60][45] = 8'h8C;
    assign wout[60][46] = 8'hC8;
    assign wout[60][47] = 8'h04;
    assign wout[60][48] = 8'h40;
    assign wout[60][49] = 8'h7C;
    assign wout[60][50] = 8'hB8;
    assign wout[60][51] = 8'hF4;
    assign wout[60][52] = 8'h30;
    assign wout[60][53] = 8'h6C;
    assign wout[60][54] = 8'hA8;
    assign wout[60][55] = 8'hE4;
    assign wout[60][56] = 8'h20;
    assign wout[60][57] = 8'h5C;
    assign wout[60][58] = 8'h98;
    assign wout[60][59] = 8'hD4;
    assign wout[60][60] = 8'h10;
    assign wout[60][61] = 8'h4C;
    assign wout[60][62] = 8'h88;
    assign wout[60][63] = 8'hC4;
    assign wout[61][0] = 8'h00;
    assign wout[61][1] = 8'h3D;
    assign wout[61][2] = 8'h7A;
    assign wout[61][3] = 8'hB7;
    assign wout[61][4] = 8'hF4;
    assign wout[61][5] = 8'h31;
    assign wout[61][6] = 8'h6E;
    assign wout[61][7] = 8'hAB;
    assign wout[61][8] = 8'hE8;
    assign wout[61][9] = 8'h25;
    assign wout[61][10] = 8'h62;
    assign wout[61][11] = 8'h9F;
    assign wout[61][12] = 8'hDC;
    assign wout[61][13] = 8'h19;
    assign wout[61][14] = 8'h56;
    assign wout[61][15] = 8'h93;
    assign wout[61][16] = 8'hD0;
    assign wout[61][17] = 8'h0D;
    assign wout[61][18] = 8'h4A;
    assign wout[61][19] = 8'h87;
    assign wout[61][20] = 8'hC4;
    assign wout[61][21] = 8'h01;
    assign wout[61][22] = 8'h3E;
    assign wout[61][23] = 8'h7B;
    assign wout[61][24] = 8'hB8;
    assign wout[61][25] = 8'hF5;
    assign wout[61][26] = 8'h32;
    assign wout[61][27] = 8'h6F;
    assign wout[61][28] = 8'hAC;
    assign wout[61][29] = 8'hE9;
    assign wout[61][30] = 8'h26;
    assign wout[61][31] = 8'h63;
    assign wout[61][32] = 8'hA0;
    assign wout[61][33] = 8'hDD;
    assign wout[61][34] = 8'h1A;
    assign wout[61][35] = 8'h57;
    assign wout[61][36] = 8'h94;
    assign wout[61][37] = 8'hD1;
    assign wout[61][38] = 8'h0E;
    assign wout[61][39] = 8'h4B;
    assign wout[61][40] = 8'h88;
    assign wout[61][41] = 8'hC5;
    assign wout[61][42] = 8'h02;
    assign wout[61][43] = 8'h3F;
    assign wout[61][44] = 8'h7C;
    assign wout[61][45] = 8'hB9;
    assign wout[61][46] = 8'hF6;
    assign wout[61][47] = 8'h33;
    assign wout[61][48] = 8'h70;
    assign wout[61][49] = 8'hAD;
    assign wout[61][50] = 8'hEA;
    assign wout[61][51] = 8'h27;
    assign wout[61][52] = 8'h64;
    assign wout[61][53] = 8'hA1;
    assign wout[61][54] = 8'hDE;
    assign wout[61][55] = 8'h1B;
    assign wout[61][56] = 8'h58;
    assign wout[61][57] = 8'h95;
    assign wout[61][58] = 8'hD2;
    assign wout[61][59] = 8'h0F;
    assign wout[61][60] = 8'h4C;
    assign wout[61][61] = 8'h89;
    assign wout[61][62] = 8'hC6;
    assign wout[61][63] = 8'h03;
    assign wout[62][0] = 8'h00;
    assign wout[62][1] = 8'h3E;
    assign wout[62][2] = 8'h7C;
    assign wout[62][3] = 8'hBA;
    assign wout[62][4] = 8'hF8;
    assign wout[62][5] = 8'h36;
    assign wout[62][6] = 8'h74;
    assign wout[62][7] = 8'hB2;
    assign wout[62][8] = 8'hF0;
    assign wout[62][9] = 8'h2E;
    assign wout[62][10] = 8'h6C;
    assign wout[62][11] = 8'hAA;
    assign wout[62][12] = 8'hE8;
    assign wout[62][13] = 8'h26;
    assign wout[62][14] = 8'h64;
    assign wout[62][15] = 8'hA2;
    assign wout[62][16] = 8'hE0;
    assign wout[62][17] = 8'h1E;
    assign wout[62][18] = 8'h5C;
    assign wout[62][19] = 8'h9A;
    assign wout[62][20] = 8'hD8;
    assign wout[62][21] = 8'h16;
    assign wout[62][22] = 8'h54;
    assign wout[62][23] = 8'h92;
    assign wout[62][24] = 8'hD0;
    assign wout[62][25] = 8'h0E;
    assign wout[62][26] = 8'h4C;
    assign wout[62][27] = 8'h8A;
    assign wout[62][28] = 8'hC8;
    assign wout[62][29] = 8'h06;
    assign wout[62][30] = 8'h44;
    assign wout[62][31] = 8'h82;
    assign wout[62][32] = 8'hC0;
    assign wout[62][33] = 8'hFE;
    assign wout[62][34] = 8'h3C;
    assign wout[62][35] = 8'h7A;
    assign wout[62][36] = 8'hB8;
    assign wout[62][37] = 8'hF6;
    assign wout[62][38] = 8'h34;
    assign wout[62][39] = 8'h72;
    assign wout[62][40] = 8'hB0;
    assign wout[62][41] = 8'hEE;
    assign wout[62][42] = 8'h2C;
    assign wout[62][43] = 8'h6A;
    assign wout[62][44] = 8'hA8;
    assign wout[62][45] = 8'hE6;
    assign wout[62][46] = 8'h24;
    assign wout[62][47] = 8'h62;
    assign wout[62][48] = 8'hA0;
    assign wout[62][49] = 8'hDE;
    assign wout[62][50] = 8'h1C;
    assign wout[62][51] = 8'h5A;
    assign wout[62][52] = 8'h98;
    assign wout[62][53] = 8'hD6;
    assign wout[62][54] = 8'h14;
    assign wout[62][55] = 8'h52;
    assign wout[62][56] = 8'h90;
    assign wout[62][57] = 8'hCE;
    assign wout[62][58] = 8'h0C;
    assign wout[62][59] = 8'h4A;
    assign wout[62][60] = 8'h88;
    assign wout[62][61] = 8'hC6;
    assign wout[62][62] = 8'h04;
    assign wout[62][63] = 8'h42;
    assign wout[63][0] = 8'h00;
    assign wout[63][1] = 8'h3F;
    assign wout[63][2] = 8'h7E;
    assign wout[63][3] = 8'hBD;
    assign wout[63][4] = 8'hFC;
    assign wout[63][5] = 8'h3B;
    assign wout[63][6] = 8'h7A;
    assign wout[63][7] = 8'hB9;
    assign wout[63][8] = 8'hF8;
    assign wout[63][9] = 8'h37;
    assign wout[63][10] = 8'h76;
    assign wout[63][11] = 8'hB5;
    assign wout[63][12] = 8'hF4;
    assign wout[63][13] = 8'h33;
    assign wout[63][14] = 8'h72;
    assign wout[63][15] = 8'hB1;
    assign wout[63][16] = 8'hF0;
    assign wout[63][17] = 8'h2F;
    assign wout[63][18] = 8'h6E;
    assign wout[63][19] = 8'hAD;
    assign wout[63][20] = 8'hEC;
    assign wout[63][21] = 8'h2B;
    assign wout[63][22] = 8'h6A;
    assign wout[63][23] = 8'hA9;
    assign wout[63][24] = 8'hE8;
    assign wout[63][25] = 8'h27;
    assign wout[63][26] = 8'h66;
    assign wout[63][27] = 8'hA5;
    assign wout[63][28] = 8'hE4;
    assign wout[63][29] = 8'h23;
    assign wout[63][30] = 8'h62;
    assign wout[63][31] = 8'hA1;
    assign wout[63][32] = 8'hE0;
    assign wout[63][33] = 8'h1F;
    assign wout[63][34] = 8'h5E;
    assign wout[63][35] = 8'h9D;
    assign wout[63][36] = 8'hDC;
    assign wout[63][37] = 8'h1B;
    assign wout[63][38] = 8'h5A;
    assign wout[63][39] = 8'h99;
    assign wout[63][40] = 8'hD8;
    assign wout[63][41] = 8'h17;
    assign wout[63][42] = 8'h56;
    assign wout[63][43] = 8'h95;
    assign wout[63][44] = 8'hD4;
    assign wout[63][45] = 8'h13;
    assign wout[63][46] = 8'h52;
    assign wout[63][47] = 8'h91;
    assign wout[63][48] = 8'hD0;
    assign wout[63][49] = 8'h0F;
    assign wout[63][50] = 8'h4E;
    assign wout[63][51] = 8'h8D;
    assign wout[63][52] = 8'hCC;
    assign wout[63][53] = 8'h0B;
    assign wout[63][54] = 8'h4A;
    assign wout[63][55] = 8'h89;
    assign wout[63][56] = 8'hC8;
    assign wout[63][57] = 8'h07;
    assign wout[63][58] = 8'h46;
    assign wout[63][59] = 8'h85;
    assign wout[63][60] = 8'hC4;
    assign wout[63][61] = 8'h03;
    assign wout[63][62] = 8'h42;
    assign wout[63][63] = 8'h81;

endmodule